`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:02:23 06/06/2015 
// Design Name: 
// Module Name:    i2s_in 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module i2s_in(
    input clk,
    input rst,
    input sck,
    input ws,
    input sd,
    output [15:0] din_lft,
    output [15:0] din_rgt,
    output din_rts,
    input din_rtr,
    output fifo_overun
    );


endmodule
