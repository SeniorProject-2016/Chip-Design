`timescale 1ns / 1ps

//////////////////////////////////////////////////////////////////////////////////
// Module Name:             reg_testbench.v
// Create Date:             2/1/2016
// Last Modification:       3/16/2016
// Author:                  Julie Swift
// Description: ????????????
//////////////////////////////////////////////////////////////////////////////////

module reg_testbench;

	// Inputs
	reg rst_n;
	reg clk;
	reg [10:0] addr;
	reg [7:0] wdata;
	reg w_enable;
	reg wxfc;
	reg ro_fifo_underrun;
	reg ro_fifo_overrun;
	reg ro_filter_ovf_flag;

	// Outputs
	wire rxfc;
	wire [7:0] rdata;
	wire rf_i2si_bist_en;
	wire [2:0] rf_filter_shift;
	wire rf_filter_clip_en;
	wire trig_fifo_overrun;
	wire trig_fifo_underrun;
	wire trig_filter_ovf_flag_clear;
	wire [7:0] rf_i2si_bist_start_val_a;
	wire [3:0] rf_i2si_bist_start_val_b;
	wire [7:0] rf_i2si_bist_incr;
	wire [7:0] rf_i2si_bist_upper_limit_a;
	wire [3:0] rf_i2si_bist_upper_limit_b;
	wire [7:0] rf_filter_coeff0_a;
	wire [7:0] rf_filter_coeff0_b;
	wire [7:0] rf_filter_coeff1_a;
	wire [7:0] rf_filter_coeff1_b;
	wire [7:0] rf_filter_coeff2_a;
	wire [7:0] rf_filter_coeff2_b;
	wire [7:0] rf_filter_coeff3_a;
	wire [7:0] rf_filter_coeff3_b;
	wire [7:0] rf_filter_coeff4_a;
	wire [7:0] rf_filter_coeff4_b;
	wire [7:0] rf_filter_coeff5_a;
	wire [7:0] rf_filter_coeff5_b;
	wire [7:0] rf_filter_coeff6_a;
	wire [7:0] rf_filter_coeff6_b;
	wire [7:0] rf_filter_coeff7_a;
	wire [7:0] rf_filter_coeff7_b;
	wire [7:0] rf_filter_coeff8_a;
	wire [7:0] rf_filter_coeff8_b;
	wire [7:0] rf_filter_coeff9_a;
	wire [7:0] rf_filter_coeff9_b;
	wire [7:0] rf_filter_coeff10_a;
	wire [7:0] rf_filter_coeff10_b;
	wire [7:0] rf_filter_coeff11_a;
	wire [7:0] rf_filter_coeff11_b;
	wire [7:0] rf_filter_coeff12_a;
	wire [7:0] rf_filter_coeff12_b;
	wire [7:0] rf_filter_coeff13_a;
	wire [7:0] rf_filter_coeff13_b;
	wire [7:0] rf_filter_coeff14_a;
	wire [7:0] rf_filter_coeff14_b;
	wire [7:0] rf_filter_coeff15_a;
	wire [7:0] rf_filter_coeff15_b;
	wire [7:0] rf_filter_coeff16_a;
	wire [7:0] rf_filter_coeff16_b;
	wire [7:0] rf_filter_coeff17_a;
	wire [7:0] rf_filter_coeff17_b;
	wire [7:0] rf_filter_coeff18_a;
	wire [7:0] rf_filter_coeff18_b;
	wire [7:0] rf_filter_coeff19_a;
	wire [7:0] rf_filter_coeff19_b;
	wire [7:0] rf_filter_coeff20_a;
	wire [7:0] rf_filter_coeff20_b;
	wire [7:0] rf_filter_coeff21_a;
	wire [7:0] rf_filter_coeff21_b;
	wire [7:0] rf_filter_coeff22_a;
	wire [7:0] rf_filter_coeff22_b;
	wire [7:0] rf_filter_coeff23_a;
	wire [7:0] rf_filter_coeff23_b;
	wire [7:0] rf_filter_coeff24_a;
	wire [7:0] rf_filter_coeff24_b;
	wire [7:0] rf_filter_coeff25_a;
	wire [7:0] rf_filter_coeff25_b;
	wire [7:0] rf_filter_coeff26_a;
	wire [7:0] rf_filter_coeff26_b;
	wire [7:0] rf_filter_coeff27_a;
	wire [7:0] rf_filter_coeff27_b;
	wire [7:0] rf_filter_coeff28_a;
	wire [7:0] rf_filter_coeff28_b;
	wire [7:0] rf_filter_coeff29_a;
	wire [7:0] rf_filter_coeff29_b;
	wire [7:0] rf_filter_coeff30_a;
	wire [7:0] rf_filter_coeff30_b;
	wire [7:0] rf_filter_coeff31_a;
	wire [7:0] rf_filter_coeff31_b;
	wire [7:0] rf_filter_coeff32_a;
	wire [7:0] rf_filter_coeff32_b;
	wire [7:0] rf_filter_coeff33_a;
	wire [7:0] rf_filter_coeff33_b;
	wire [7:0] rf_filter_coeff34_a;
	wire [7:0] rf_filter_coeff34_b;
	wire [7:0] rf_filter_coeff35_a;
	wire [7:0] rf_filter_coeff35_b;
	wire [7:0] rf_filter_coeff36_a;
	wire [7:0] rf_filter_coeff36_b;
	wire [7:0] rf_filter_coeff37_a;
	wire [7:0] rf_filter_coeff37_b;
	wire [7:0] rf_filter_coeff38_a;
	wire [7:0] rf_filter_coeff38_b;
	wire [7:0] rf_filter_coeff39_a;
	wire [7:0] rf_filter_coeff39_b;
	wire [7:0] rf_filter_coeff40_a;
	wire [7:0] rf_filter_coeff40_b;
	wire [7:0] rf_filter_coeff41_a;
	wire [7:0] rf_filter_coeff41_b;
	wire [7:0] rf_filter_coeff42_a;
	wire [7:0] rf_filter_coeff42_b;
	wire [7:0] rf_filter_coeff43_a;
	wire [7:0] rf_filter_coeff43_b;
	wire [7:0] rf_filter_coeff44_a;
	wire [7:0] rf_filter_coeff44_b;
	wire [7:0] rf_filter_coeff45_a;
	wire [7:0] rf_filter_coeff45_b;
	wire [7:0] rf_filter_coeff46_a;
	wire [7:0] rf_filter_coeff46_b;
	wire [7:0] rf_filter_coeff47_a;
	wire [7:0] rf_filter_coeff47_b;
	wire [7:0] rf_filter_coeff48_a;
	wire [7:0] rf_filter_coeff48_b;
	wire [7:0] rf_filter_coeff49_a;
	wire [7:0] rf_filter_coeff49_b;
	wire [7:0] rf_filter_coeff50_a;
	wire [7:0] rf_filter_coeff50_b;
	wire [7:0] rf_filter_coeff51_a;
	wire [7:0] rf_filter_coeff51_b;
	wire [7:0] rf_filter_coeff52_a;
	wire [7:0] rf_filter_coeff52_b;
	wire [7:0] rf_filter_coeff53_a;
	wire [7:0] rf_filter_coeff53_b;
	wire [7:0] rf_filter_coeff54_a;
	wire [7:0] rf_filter_coeff54_b;
	wire [7:0] rf_filter_coeff55_a;
	wire [7:0] rf_filter_coeff55_b;
	wire [7:0] rf_filter_coeff56_a;
	wire [7:0] rf_filter_coeff56_b;
	wire [7:0] rf_filter_coeff57_a;
	wire [7:0] rf_filter_coeff57_b;
	wire [7:0] rf_filter_coeff58_a;
	wire [7:0] rf_filter_coeff58_b;
	wire [7:0] rf_filter_coeff59_a;
	wire [7:0] rf_filter_coeff59_b;
	wire [7:0] rf_filter_coeff60_a;
	wire [7:0] rf_filter_coeff60_b;
	wire [7:0] rf_filter_coeff61_a;
	wire [7:0] rf_filter_coeff61_b;
	wire [7:0] rf_filter_coeff62_a;
	wire [7:0] rf_filter_coeff62_b;
	wire [7:0] rf_filter_coeff63_a;
	wire [7:0] rf_filter_coeff63_b;
	wire [7:0] rf_filter_coeff64_a;
	wire [7:0] rf_filter_coeff64_b;
	wire [7:0] rf_filter_coeff65_a;
	wire [7:0] rf_filter_coeff65_b;
	wire [7:0] rf_filter_coeff66_a;
	wire [7:0] rf_filter_coeff66_b;
	wire [7:0] rf_filter_coeff67_a;
	wire [7:0] rf_filter_coeff67_b;
	wire [7:0] rf_filter_coeff68_a;
	wire [7:0] rf_filter_coeff68_b;
	wire [7:0] rf_filter_coeff69_a;
	wire [7:0] rf_filter_coeff69_b;
	wire [7:0] rf_filter_coeff70_a;
	wire [7:0] rf_filter_coeff70_b;
	wire [7:0] rf_filter_coeff71_a;
	wire [7:0] rf_filter_coeff71_b;
	wire [7:0] rf_filter_coeff72_a;
	wire [7:0] rf_filter_coeff72_b;
	wire [7:0] rf_filter_coeff73_a;
	wire [7:0] rf_filter_coeff73_b;
	wire [7:0] rf_filter_coeff74_a;
	wire [7:0] rf_filter_coeff74_b;
	wire [7:0] rf_filter_coeff75_a;
	wire [7:0] rf_filter_coeff75_b;
	wire [7:0] rf_filter_coeff76_a;
	wire [7:0] rf_filter_coeff76_b;
	wire [7:0] rf_filter_coeff77_a;
	wire [7:0] rf_filter_coeff77_b;
	wire [7:0] rf_filter_coeff78_a;
	wire [7:0] rf_filter_coeff78_b;
	wire [7:0] rf_filter_coeff79_a;
	wire [7:0] rf_filter_coeff79_b;
	wire [7:0] rf_filter_coeff80_a;
	wire [7:0] rf_filter_coeff80_b;
	wire [7:0] rf_filter_coeff81_a;
	wire [7:0] rf_filter_coeff81_b;
	wire [7:0] rf_filter_coeff82_a;
	wire [7:0] rf_filter_coeff82_b;
	wire [7:0] rf_filter_coeff83_a;
	wire [7:0] rf_filter_coeff83_b;
	wire [7:0] rf_filter_coeff84_a;
	wire [7:0] rf_filter_coeff84_b;
	wire [7:0] rf_filter_coeff85_a;
	wire [7:0] rf_filter_coeff85_b;
	wire [7:0] rf_filter_coeff86_a;
	wire [7:0] rf_filter_coeff86_b;
	wire [7:0] rf_filter_coeff87_a;
	wire [7:0] rf_filter_coeff87_b;
	wire [7:0] rf_filter_coeff88_a;
	wire [7:0] rf_filter_coeff88_b;
	wire [7:0] rf_filter_coeff89_a;
	wire [7:0] rf_filter_coeff89_b;
	wire [7:0] rf_filter_coeff90_a;
	wire [7:0] rf_filter_coeff90_b;
	wire [7:0] rf_filter_coeff91_a;
	wire [7:0] rf_filter_coeff91_b;
	wire [7:0] rf_filter_coeff92_a;
	wire [7:0] rf_filter_coeff92_b;
	wire [7:0] rf_filter_coeff93_a;
	wire [7:0] rf_filter_coeff93_b;
	wire [7:0] rf_filter_coeff94_a;
	wire [7:0] rf_filter_coeff94_b;
	wire [7:0] rf_filter_coeff95_a;
	wire [7:0] rf_filter_coeff95_b;
	wire [7:0] rf_filter_coeff96_a;
	wire [7:0] rf_filter_coeff96_b;
	wire [7:0] rf_filter_coeff97_a;
	wire [7:0] rf_filter_coeff97_b;
	wire [7:0] rf_filter_coeff98_a;
	wire [7:0] rf_filter_coeff98_b;
	wire [7:0] rf_filter_coeff99_a;
	wire [7:0] rf_filter_coeff99_b;
	wire [7:0] rf_filter_coeff100_a;
	wire [7:0] rf_filter_coeff100_b;
	wire [7:0] rf_filter_coeff101_a;
	wire [7:0] rf_filter_coeff101_b;
	wire [7:0] rf_filter_coeff102_a;
	wire [7:0] rf_filter_coeff102_b;
	wire [7:0] rf_filter_coeff103_a;
	wire [7:0] rf_filter_coeff103_b;
	wire [7:0] rf_filter_coeff104_a;
	wire [7:0] rf_filter_coeff104_b;
	wire [7:0] rf_filter_coeff105_a;
	wire [7:0] rf_filter_coeff105_b;
	wire [7:0] rf_filter_coeff106_a;
	wire [7:0] rf_filter_coeff106_b;
	wire [7:0] rf_filter_coeff107_a;
	wire [7:0] rf_filter_coeff107_b;
	wire [7:0] rf_filter_coeff108_a;
	wire [7:0] rf_filter_coeff108_b;
	wire [7:0] rf_filter_coeff109_a;
	wire [7:0] rf_filter_coeff109_b;
	wire [7:0] rf_filter_coeff110_a;
	wire [7:0] rf_filter_coeff110_b;
	wire [7:0] rf_filter_coeff111_a;
	wire [7:0] rf_filter_coeff111_b;
	wire [7:0] rf_filter_coeff112_a;
	wire [7:0] rf_filter_coeff112_b;
	wire [7:0] rf_filter_coeff113_a;
	wire [7:0] rf_filter_coeff113_b;
	wire [7:0] rf_filter_coeff114_a;
	wire [7:0] rf_filter_coeff114_b;
	wire [7:0] rf_filter_coeff115_a;
	wire [7:0] rf_filter_coeff115_b;
	wire [7:0] rf_filter_coeff116_a;
	wire [7:0] rf_filter_coeff116_b;
	wire [7:0] rf_filter_coeff117_a;
	wire [7:0] rf_filter_coeff117_b;
	wire [7:0] rf_filter_coeff118_a;
	wire [7:0] rf_filter_coeff118_b;
	wire [7:0] rf_filter_coeff119_a;
	wire [7:0] rf_filter_coeff119_b;
	wire [7:0] rf_filter_coeff120_a;
	wire [7:0] rf_filter_coeff120_b;
	wire [7:0] rf_filter_coeff121_a;
	wire [7:0] rf_filter_coeff121_b;
	wire [7:0] rf_filter_coeff122_a;
	wire [7:0] rf_filter_coeff122_b;
	wire [7:0] rf_filter_coeff123_a;
	wire [7:0] rf_filter_coeff123_b;
	wire [7:0] rf_filter_coeff124_a;
	wire [7:0] rf_filter_coeff124_b;
	wire [7:0] rf_filter_coeff125_a;
	wire [7:0] rf_filter_coeff125_b;
	wire [7:0] rf_filter_coeff126_a;
	wire [7:0] rf_filter_coeff126_b;
	wire [7:0] rf_filter_coeff127_a;
	wire [7:0] rf_filter_coeff127_b;
	wire [7:0] rf_filter_coeff128_a;
	wire [7:0] rf_filter_coeff128_b;
	wire [7:0] rf_filter_coeff129_a;
	wire [7:0] rf_filter_coeff129_b;
	wire [7:0] rf_filter_coeff130_a;
	wire [7:0] rf_filter_coeff130_b;
	wire [7:0] rf_filter_coeff131_a;
	wire [7:0] rf_filter_coeff131_b;
	wire [7:0] rf_filter_coeff132_a;
	wire [7:0] rf_filter_coeff132_b;
	wire [7:0] rf_filter_coeff133_a;
	wire [7:0] rf_filter_coeff133_b;
	wire [7:0] rf_filter_coeff134_a;
	wire [7:0] rf_filter_coeff134_b;
	wire [7:0] rf_filter_coeff135_a;
	wire [7:0] rf_filter_coeff135_b;
	wire [7:0] rf_filter_coeff136_a;
	wire [7:0] rf_filter_coeff136_b;
	wire [7:0] rf_filter_coeff137_a;
	wire [7:0] rf_filter_coeff137_b;
	wire [7:0] rf_filter_coeff138_a;
	wire [7:0] rf_filter_coeff138_b;
	wire [7:0] rf_filter_coeff139_a;
	wire [7:0] rf_filter_coeff139_b;
	wire [7:0] rf_filter_coeff140_a;
	wire [7:0] rf_filter_coeff140_b;
	wire [7:0] rf_filter_coeff141_a;
	wire [7:0] rf_filter_coeff141_b;
	wire [7:0] rf_filter_coeff142_a;
	wire [7:0] rf_filter_coeff142_b;
	wire [7:0] rf_filter_coeff143_a;
	wire [7:0] rf_filter_coeff143_b;
	wire [7:0] rf_filter_coeff144_a;
	wire [7:0] rf_filter_coeff144_b;
	wire [7:0] rf_filter_coeff145_a;
	wire [7:0] rf_filter_coeff145_b;
	wire [7:0] rf_filter_coeff146_a;
	wire [7:0] rf_filter_coeff146_b;
	wire [7:0] rf_filter_coeff147_a;
	wire [7:0] rf_filter_coeff147_b;
	wire [7:0] rf_filter_coeff148_a;
	wire [7:0] rf_filter_coeff148_b;
	wire [7:0] rf_filter_coeff149_a;
	wire [7:0] rf_filter_coeff149_b;
	wire [7:0] rf_filter_coeff150_a;
	wire [7:0] rf_filter_coeff150_b;
	wire [7:0] rf_filter_coeff151_a;
	wire [7:0] rf_filter_coeff151_b;
	wire [7:0] rf_filter_coeff152_a;
	wire [7:0] rf_filter_coeff152_b;
	wire [7:0] rf_filter_coeff153_a;
	wire [7:0] rf_filter_coeff153_b;
	wire [7:0] rf_filter_coeff154_a;
	wire [7:0] rf_filter_coeff154_b;
	wire [7:0] rf_filter_coeff155_a;
	wire [7:0] rf_filter_coeff155_b;
	wire [7:0] rf_filter_coeff156_a;
	wire [7:0] rf_filter_coeff156_b;
	wire [7:0] rf_filter_coeff157_a;
	wire [7:0] rf_filter_coeff157_b;
	wire [7:0] rf_filter_coeff158_a;
	wire [7:0] rf_filter_coeff158_b;
	wire [7:0] rf_filter_coeff159_a;
	wire [7:0] rf_filter_coeff159_b;
	wire [7:0] rf_filter_coeff160_a;
	wire [7:0] rf_filter_coeff160_b;
	wire [7:0] rf_filter_coeff161_a;
	wire [7:0] rf_filter_coeff161_b;
	wire [7:0] rf_filter_coeff162_a;
	wire [7:0] rf_filter_coeff162_b;
	wire [7:0] rf_filter_coeff163_a;
	wire [7:0] rf_filter_coeff163_b;
	wire [7:0] rf_filter_coeff164_a;
	wire [7:0] rf_filter_coeff164_b;
	wire [7:0] rf_filter_coeff165_a;
	wire [7:0] rf_filter_coeff165_b;
	wire [7:0] rf_filter_coeff166_a;
	wire [7:0] rf_filter_coeff166_b;
	wire [7:0] rf_filter_coeff167_a;
	wire [7:0] rf_filter_coeff167_b;
	wire [7:0] rf_filter_coeff168_a;
	wire [7:0] rf_filter_coeff168_b;
	wire [7:0] rf_filter_coeff169_a;
	wire [7:0] rf_filter_coeff169_b;
	wire [7:0] rf_filter_coeff170_a;
	wire [7:0] rf_filter_coeff170_b;
	wire [7:0] rf_filter_coeff171_a;
	wire [7:0] rf_filter_coeff171_b;
	wire [7:0] rf_filter_coeff172_a;
	wire [7:0] rf_filter_coeff172_b;
	wire [7:0] rf_filter_coeff173_a;
	wire [7:0] rf_filter_coeff173_b;
	wire [7:0] rf_filter_coeff174_a;
	wire [7:0] rf_filter_coeff174_b;
	wire [7:0] rf_filter_coeff175_a;
	wire [7:0] rf_filter_coeff175_b;
	wire [7:0] rf_filter_coeff176_a;
	wire [7:0] rf_filter_coeff176_b;
	wire [7:0] rf_filter_coeff177_a;
	wire [7:0] rf_filter_coeff177_b;
	wire [7:0] rf_filter_coeff178_a;
	wire [7:0] rf_filter_coeff178_b;
	wire [7:0] rf_filter_coeff179_a;
	wire [7:0] rf_filter_coeff179_b;
	wire [7:0] rf_filter_coeff180_a;
	wire [7:0] rf_filter_coeff180_b;
	wire [7:0] rf_filter_coeff181_a;
	wire [7:0] rf_filter_coeff181_b;
	wire [7:0] rf_filter_coeff182_a;
	wire [7:0] rf_filter_coeff182_b;
	wire [7:0] rf_filter_coeff183_a;
	wire [7:0] rf_filter_coeff183_b;
	wire [7:0] rf_filter_coeff184_a;
	wire [7:0] rf_filter_coeff184_b;
	wire [7:0] rf_filter_coeff185_a;
	wire [7:0] rf_filter_coeff185_b;
	wire [7:0] rf_filter_coeff186_a;
	wire [7:0] rf_filter_coeff186_b;
	wire [7:0] rf_filter_coeff187_a;
	wire [7:0] rf_filter_coeff187_b;
	wire [7:0] rf_filter_coeff188_a;
	wire [7:0] rf_filter_coeff188_b;
	wire [7:0] rf_filter_coeff189_a;
	wire [7:0] rf_filter_coeff189_b;
	wire [7:0] rf_filter_coeff190_a;
	wire [7:0] rf_filter_coeff190_b;
	wire [7:0] rf_filter_coeff191_a;
	wire [7:0] rf_filter_coeff191_b;
	wire [7:0] rf_filter_coeff192_a;
	wire [7:0] rf_filter_coeff192_b;
	wire [7:0] rf_filter_coeff193_a;
	wire [7:0] rf_filter_coeff193_b;
	wire [7:0] rf_filter_coeff194_a;
	wire [7:0] rf_filter_coeff194_b;
	wire [7:0] rf_filter_coeff195_a;
	wire [7:0] rf_filter_coeff195_b;
	wire [7:0] rf_filter_coeff196_a;
	wire [7:0] rf_filter_coeff196_b;
	wire [7:0] rf_filter_coeff197_a;
	wire [7:0] rf_filter_coeff197_b;
	wire [7:0] rf_filter_coeff198_a;
	wire [7:0] rf_filter_coeff198_b;
	wire [7:0] rf_filter_coeff199_a;
	wire [7:0] rf_filter_coeff199_b;
	wire [7:0] rf_filter_coeff200_a;
	wire [7:0] rf_filter_coeff200_b;
	wire [7:0] rf_filter_coeff201_a;
	wire [7:0] rf_filter_coeff201_b;
	wire [7:0] rf_filter_coeff202_a;
	wire [7:0] rf_filter_coeff202_b;
	wire [7:0] rf_filter_coeff203_a;
	wire [7:0] rf_filter_coeff203_b;
	wire [7:0] rf_filter_coeff204_a;
	wire [7:0] rf_filter_coeff204_b;
	wire [7:0] rf_filter_coeff205_a;
	wire [7:0] rf_filter_coeff205_b;
	wire [7:0] rf_filter_coeff206_a;
	wire [7:0] rf_filter_coeff206_b;
	wire [7:0] rf_filter_coeff207_a;
	wire [7:0] rf_filter_coeff207_b;
	wire [7:0] rf_filter_coeff208_a;
	wire [7:0] rf_filter_coeff208_b;
	wire [7:0] rf_filter_coeff209_a;
	wire [7:0] rf_filter_coeff209_b;
	wire [7:0] rf_filter_coeff210_a;
	wire [7:0] rf_filter_coeff210_b;
	wire [7:0] rf_filter_coeff211_a;
	wire [7:0] rf_filter_coeff211_b;
	wire [7:0] rf_filter_coeff212_a;
	wire [7:0] rf_filter_coeff212_b;
	wire [7:0] rf_filter_coeff213_a;
	wire [7:0] rf_filter_coeff213_b;
	wire [7:0] rf_filter_coeff214_a;
	wire [7:0] rf_filter_coeff214_b;
	wire [7:0] rf_filter_coeff215_a;
	wire [7:0] rf_filter_coeff215_b;
	wire [7:0] rf_filter_coeff216_a;
	wire [7:0] rf_filter_coeff216_b;
	wire [7:0] rf_filter_coeff217_a;
	wire [7:0] rf_filter_coeff217_b;
	wire [7:0] rf_filter_coeff218_a;
	wire [7:0] rf_filter_coeff218_b;
	wire [7:0] rf_filter_coeff219_a;
	wire [7:0] rf_filter_coeff219_b;
	wire [7:0] rf_filter_coeff220_a;
	wire [7:0] rf_filter_coeff220_b;
	wire [7:0] rf_filter_coeff221_a;
	wire [7:0] rf_filter_coeff221_b;
	wire [7:0] rf_filter_coeff222_a;
	wire [7:0] rf_filter_coeff222_b;
	wire [7:0] rf_filter_coeff223_a;
	wire [7:0] rf_filter_coeff223_b;
	wire [7:0] rf_filter_coeff224_a;
	wire [7:0] rf_filter_coeff224_b;
	wire [7:0] rf_filter_coeff225_a;
	wire [7:0] rf_filter_coeff225_b;
	wire [7:0] rf_filter_coeff226_a;
	wire [7:0] rf_filter_coeff226_b;
	wire [7:0] rf_filter_coeff227_a;
	wire [7:0] rf_filter_coeff227_b;
	wire [7:0] rf_filter_coeff228_a;
	wire [7:0] rf_filter_coeff228_b;
	wire [7:0] rf_filter_coeff229_a;
	wire [7:0] rf_filter_coeff229_b;
	wire [7:0] rf_filter_coeff230_a;
	wire [7:0] rf_filter_coeff230_b;
	wire [7:0] rf_filter_coeff231_a;
	wire [7:0] rf_filter_coeff231_b;
	wire [7:0] rf_filter_coeff232_a;
	wire [7:0] rf_filter_coeff232_b;
	wire [7:0] rf_filter_coeff233_a;
	wire [7:0] rf_filter_coeff233_b;
	wire [7:0] rf_filter_coeff234_a;
	wire [7:0] rf_filter_coeff234_b;
	wire [7:0] rf_filter_coeff235_a;
	wire [7:0] rf_filter_coeff235_b;
	wire [7:0] rf_filter_coeff236_a;
	wire [7:0] rf_filter_coeff236_b;
	wire [7:0] rf_filter_coeff237_a;
	wire [7:0] rf_filter_coeff237_b;
	wire [7:0] rf_filter_coeff238_a;
	wire [7:0] rf_filter_coeff238_b;
	wire [7:0] rf_filter_coeff239_a;
	wire [7:0] rf_filter_coeff239_b;
	wire [7:0] rf_filter_coeff240_a;
	wire [7:0] rf_filter_coeff240_b;
	wire [7:0] rf_filter_coeff241_a;
	wire [7:0] rf_filter_coeff241_b;
	wire [7:0] rf_filter_coeff242_a;
	wire [7:0] rf_filter_coeff242_b;
	wire [7:0] rf_filter_coeff243_a;
	wire [7:0] rf_filter_coeff243_b;
	wire [7:0] rf_filter_coeff244_a;
	wire [7:0] rf_filter_coeff244_b;
	wire [7:0] rf_filter_coeff245_a;
	wire [7:0] rf_filter_coeff245_b;
	wire [7:0] rf_filter_coeff246_a;
	wire [7:0] rf_filter_coeff246_b;
	wire [7:0] rf_filter_coeff247_a;
	wire [7:0] rf_filter_coeff247_b;
	wire [7:0] rf_filter_coeff248_a;
	wire [7:0] rf_filter_coeff248_b;
	wire [7:0] rf_filter_coeff249_a;
	wire [7:0] rf_filter_coeff249_b;
	wire [7:0] rf_filter_coeff250_a;
	wire [7:0] rf_filter_coeff250_b;
	wire [7:0] rf_filter_coeff251_a;
	wire [7:0] rf_filter_coeff251_b;
	wire [7:0] rf_filter_coeff252_a;
	wire [7:0] rf_filter_coeff252_b;
	wire [7:0] rf_filter_coeff253_a;
	wire [7:0] rf_filter_coeff253_b;
	wire [7:0] rf_filter_coeff254_a;
	wire [7:0] rf_filter_coeff254_b;
	wire [7:0] rf_filter_coeff255_a;
	wire [7:0] rf_filter_coeff255_b;
	wire [7:0] rf_filter_coeff256_a;
	wire [7:0] rf_filter_coeff256_b;
	wire [7:0] rf_filter_coeff257_a;
	wire [7:0] rf_filter_coeff257_b;
	wire [7:0] rf_filter_coeff258_a;
	wire [7:0] rf_filter_coeff258_b;
	wire [7:0] rf_filter_coeff259_a;
	wire [7:0] rf_filter_coeff259_b;
	wire [7:0] rf_filter_coeff260_a;
	wire [7:0] rf_filter_coeff260_b;
	wire [7:0] rf_filter_coeff261_a;
	wire [7:0] rf_filter_coeff261_b;
	wire [7:0] rf_filter_coeff262_a;
	wire [7:0] rf_filter_coeff262_b;
	wire [7:0] rf_filter_coeff263_a;
	wire [7:0] rf_filter_coeff263_b;
	wire [7:0] rf_filter_coeff264_a;
	wire [7:0] rf_filter_coeff264_b;
	wire [7:0] rf_filter_coeff265_a;
	wire [7:0] rf_filter_coeff265_b;
	wire [7:0] rf_filter_coeff266_a;
	wire [7:0] rf_filter_coeff266_b;
	wire [7:0] rf_filter_coeff267_a;
	wire [7:0] rf_filter_coeff267_b;
	wire [7:0] rf_filter_coeff268_a;
	wire [7:0] rf_filter_coeff268_b;
	wire [7:0] rf_filter_coeff269_a;
	wire [7:0] rf_filter_coeff269_b;
	wire [7:0] rf_filter_coeff270_a;
	wire [7:0] rf_filter_coeff270_b;
	wire [7:0] rf_filter_coeff271_a;
	wire [7:0] rf_filter_coeff271_b;
	wire [7:0] rf_filter_coeff272_a;
	wire [7:0] rf_filter_coeff272_b;
	wire [7:0] rf_filter_coeff273_a;
	wire [7:0] rf_filter_coeff273_b;
	wire [7:0] rf_filter_coeff274_a;
	wire [7:0] rf_filter_coeff274_b;
	wire [7:0] rf_filter_coeff275_a;
	wire [7:0] rf_filter_coeff275_b;
	wire [7:0] rf_filter_coeff276_a;
	wire [7:0] rf_filter_coeff276_b;
	wire [7:0] rf_filter_coeff277_a;
	wire [7:0] rf_filter_coeff277_b;
	wire [7:0] rf_filter_coeff278_a;
	wire [7:0] rf_filter_coeff278_b;
	wire [7:0] rf_filter_coeff279_a;
	wire [7:0] rf_filter_coeff279_b;
	wire [7:0] rf_filter_coeff280_a;
	wire [7:0] rf_filter_coeff280_b;
	wire [7:0] rf_filter_coeff281_a;
	wire [7:0] rf_filter_coeff281_b;
	wire [7:0] rf_filter_coeff282_a;
	wire [7:0] rf_filter_coeff282_b;
	wire [7:0] rf_filter_coeff283_a;
	wire [7:0] rf_filter_coeff283_b;
	wire [7:0] rf_filter_coeff284_a;
	wire [7:0] rf_filter_coeff284_b;
	wire [7:0] rf_filter_coeff285_a;
	wire [7:0] rf_filter_coeff285_b;
	wire [7:0] rf_filter_coeff286_a;
	wire [7:0] rf_filter_coeff286_b;
	wire [7:0] rf_filter_coeff287_a;
	wire [7:0] rf_filter_coeff287_b;
	wire [7:0] rf_filter_coeff288_a;
	wire [7:0] rf_filter_coeff288_b;
	wire [7:0] rf_filter_coeff289_a;
	wire [7:0] rf_filter_coeff289_b;
	wire [7:0] rf_filter_coeff290_a;
	wire [7:0] rf_filter_coeff290_b;
	wire [7:0] rf_filter_coeff291_a;
	wire [7:0] rf_filter_coeff291_b;
	wire [7:0] rf_filter_coeff292_a;
	wire [7:0] rf_filter_coeff292_b;
	wire [7:0] rf_filter_coeff293_a;
	wire [7:0] rf_filter_coeff293_b;
	wire [7:0] rf_filter_coeff294_a;
	wire [7:0] rf_filter_coeff294_b;
	wire [7:0] rf_filter_coeff295_a;
	wire [7:0] rf_filter_coeff295_b;
	wire [7:0] rf_filter_coeff296_a;
	wire [7:0] rf_filter_coeff296_b;
	wire [7:0] rf_filter_coeff297_a;
	wire [7:0] rf_filter_coeff297_b;
	wire [7:0] rf_filter_coeff298_a;
	wire [7:0] rf_filter_coeff298_b;
	wire [7:0] rf_filter_coeff299_a;
	wire [7:0] rf_filter_coeff299_b;
	wire [7:0] rf_filter_coeff300_a;
	wire [7:0] rf_filter_coeff300_b;
	wire [7:0] rf_filter_coeff301_a;
	wire [7:0] rf_filter_coeff301_b;
	wire [7:0] rf_filter_coeff302_a;
	wire [7:0] rf_filter_coeff302_b;
	wire [7:0] rf_filter_coeff303_a;
	wire [7:0] rf_filter_coeff303_b;
	wire [7:0] rf_filter_coeff304_a;
	wire [7:0] rf_filter_coeff304_b;
	wire [7:0] rf_filter_coeff305_a;
	wire [7:0] rf_filter_coeff305_b;
	wire [7:0] rf_filter_coeff306_a;
	wire [7:0] rf_filter_coeff306_b;
	wire [7:0] rf_filter_coeff307_a;
	wire [7:0] rf_filter_coeff307_b;
	wire [7:0] rf_filter_coeff308_a;
	wire [7:0] rf_filter_coeff308_b;
	wire [7:0] rf_filter_coeff309_a;
	wire [7:0] rf_filter_coeff309_b;
	wire [7:0] rf_filter_coeff310_a;
	wire [7:0] rf_filter_coeff310_b;
	wire [7:0] rf_filter_coeff311_a;
	wire [7:0] rf_filter_coeff311_b;
	wire [7:0] rf_filter_coeff312_a;
	wire [7:0] rf_filter_coeff312_b;
	wire [7:0] rf_filter_coeff313_a;
	wire [7:0] rf_filter_coeff313_b;
	wire [7:0] rf_filter_coeff314_a;
	wire [7:0] rf_filter_coeff314_b;
	wire [7:0] rf_filter_coeff315_a;
	wire [7:0] rf_filter_coeff315_b;
	wire [7:0] rf_filter_coeff316_a;
	wire [7:0] rf_filter_coeff316_b;
	wire [7:0] rf_filter_coeff317_a;
	wire [7:0] rf_filter_coeff317_b;
	wire [7:0] rf_filter_coeff318_a;
	wire [7:0] rf_filter_coeff318_b;
	wire [7:0] rf_filter_coeff319_a;
	wire [7:0] rf_filter_coeff319_b;
	wire [7:0] rf_filter_coeff320_a;
	wire [7:0] rf_filter_coeff320_b;
	wire [7:0] rf_filter_coeff321_a;
	wire [7:0] rf_filter_coeff321_b;
	wire [7:0] rf_filter_coeff322_a;
	wire [7:0] rf_filter_coeff322_b;
	wire [7:0] rf_filter_coeff323_a;
	wire [7:0] rf_filter_coeff323_b;
	wire [7:0] rf_filter_coeff324_a;
	wire [7:0] rf_filter_coeff324_b;
	wire [7:0] rf_filter_coeff325_a;
	wire [7:0] rf_filter_coeff325_b;
	wire [7:0] rf_filter_coeff326_a;
	wire [7:0] rf_filter_coeff326_b;
	wire [7:0] rf_filter_coeff327_a;
	wire [7:0] rf_filter_coeff327_b;
	wire [7:0] rf_filter_coeff328_a;
	wire [7:0] rf_filter_coeff328_b;
	wire [7:0] rf_filter_coeff329_a;
	wire [7:0] rf_filter_coeff329_b;
	wire [7:0] rf_filter_coeff330_a;
	wire [7:0] rf_filter_coeff330_b;
	wire [7:0] rf_filter_coeff331_a;
	wire [7:0] rf_filter_coeff331_b;
	wire [7:0] rf_filter_coeff332_a;
	wire [7:0] rf_filter_coeff332_b;
	wire [7:0] rf_filter_coeff333_a;
	wire [7:0] rf_filter_coeff333_b;
	wire [7:0] rf_filter_coeff334_a;
	wire [7:0] rf_filter_coeff334_b;
	wire [7:0] rf_filter_coeff335_a;
	wire [7:0] rf_filter_coeff335_b;
	wire [7:0] rf_filter_coeff336_a;
	wire [7:0] rf_filter_coeff336_b;
	wire [7:0] rf_filter_coeff337_a;
	wire [7:0] rf_filter_coeff337_b;
	wire [7:0] rf_filter_coeff338_a;
	wire [7:0] rf_filter_coeff338_b;
	wire [7:0] rf_filter_coeff339_a;
	wire [7:0] rf_filter_coeff339_b;
	wire [7:0] rf_filter_coeff340_a;
	wire [7:0] rf_filter_coeff340_b;
	wire [7:0] rf_filter_coeff341_a;
	wire [7:0] rf_filter_coeff341_b;
	wire [7:0] rf_filter_coeff342_a;
	wire [7:0] rf_filter_coeff342_b;
	wire [7:0] rf_filter_coeff343_a;
	wire [7:0] rf_filter_coeff343_b;
	wire [7:0] rf_filter_coeff344_a;
	wire [7:0] rf_filter_coeff344_b;
	wire [7:0] rf_filter_coeff345_a;
	wire [7:0] rf_filter_coeff345_b;
	wire [7:0] rf_filter_coeff346_a;
	wire [7:0] rf_filter_coeff346_b;
	wire [7:0] rf_filter_coeff347_a;
	wire [7:0] rf_filter_coeff347_b;
	wire [7:0] rf_filter_coeff348_a;
	wire [7:0] rf_filter_coeff348_b;
	wire [7:0] rf_filter_coeff349_a;
	wire [7:0] rf_filter_coeff349_b;
	wire [7:0] rf_filter_coeff350_a;
	wire [7:0] rf_filter_coeff350_b;
	wire [7:0] rf_filter_coeff351_a;
	wire [7:0] rf_filter_coeff351_b;
	wire [7:0] rf_filter_coeff352_a;
	wire [7:0] rf_filter_coeff352_b;
	wire [7:0] rf_filter_coeff353_a;
	wire [7:0] rf_filter_coeff353_b;
	wire [7:0] rf_filter_coeff354_a;
	wire [7:0] rf_filter_coeff354_b;
	wire [7:0] rf_filter_coeff355_a;
	wire [7:0] rf_filter_coeff355_b;
	wire [7:0] rf_filter_coeff356_a;
	wire [7:0] rf_filter_coeff356_b;
	wire [7:0] rf_filter_coeff357_a;
	wire [7:0] rf_filter_coeff357_b;
	wire [7:0] rf_filter_coeff358_a;
	wire [7:0] rf_filter_coeff358_b;
	wire [7:0] rf_filter_coeff359_a;
	wire [7:0] rf_filter_coeff359_b;
	wire [7:0] rf_filter_coeff360_a;
	wire [7:0] rf_filter_coeff360_b;
	wire [7:0] rf_filter_coeff361_a;
	wire [7:0] rf_filter_coeff361_b;
	wire [7:0] rf_filter_coeff362_a;
	wire [7:0] rf_filter_coeff362_b;
	wire [7:0] rf_filter_coeff363_a;
	wire [7:0] rf_filter_coeff363_b;
	wire [7:0] rf_filter_coeff364_a;
	wire [7:0] rf_filter_coeff364_b;
	wire [7:0] rf_filter_coeff365_a;
	wire [7:0] rf_filter_coeff365_b;
	wire [7:0] rf_filter_coeff366_a;
	wire [7:0] rf_filter_coeff366_b;
	wire [7:0] rf_filter_coeff367_a;
	wire [7:0] rf_filter_coeff367_b;
	wire [7:0] rf_filter_coeff368_a;
	wire [7:0] rf_filter_coeff368_b;
	wire [7:0] rf_filter_coeff369_a;
	wire [7:0] rf_filter_coeff369_b;
	wire [7:0] rf_filter_coeff370_a;
	wire [7:0] rf_filter_coeff370_b;
	wire [7:0] rf_filter_coeff371_a;
	wire [7:0] rf_filter_coeff371_b;
	wire [7:0] rf_filter_coeff372_a;
	wire [7:0] rf_filter_coeff372_b;
	wire [7:0] rf_filter_coeff373_a;
	wire [7:0] rf_filter_coeff373_b;
	wire [7:0] rf_filter_coeff374_a;
	wire [7:0] rf_filter_coeff374_b;
	wire [7:0] rf_filter_coeff375_a;
	wire [7:0] rf_filter_coeff375_b;
	wire [7:0] rf_filter_coeff376_a;
	wire [7:0] rf_filter_coeff376_b;
	wire [7:0] rf_filter_coeff377_a;
	wire [7:0] rf_filter_coeff377_b;
	wire [7:0] rf_filter_coeff378_a;
	wire [7:0] rf_filter_coeff378_b;
	wire [7:0] rf_filter_coeff379_a;
	wire [7:0] rf_filter_coeff379_b;
	wire [7:0] rf_filter_coeff380_a;
	wire [7:0] rf_filter_coeff380_b;
	wire [7:0] rf_filter_coeff381_a;
	wire [7:0] rf_filter_coeff381_b;
	wire [7:0] rf_filter_coeff382_a;
	wire [7:0] rf_filter_coeff382_b;
	wire [7:0] rf_filter_coeff383_a;
	wire [7:0] rf_filter_coeff383_b;
	wire [7:0] rf_filter_coeff384_a;
	wire [7:0] rf_filter_coeff384_b;
	wire [7:0] rf_filter_coeff385_a;
	wire [7:0] rf_filter_coeff385_b;
	wire [7:0] rf_filter_coeff386_a;
	wire [7:0] rf_filter_coeff386_b;
	wire [7:0] rf_filter_coeff387_a;
	wire [7:0] rf_filter_coeff387_b;
	wire [7:0] rf_filter_coeff388_a;
	wire [7:0] rf_filter_coeff388_b;
	wire [7:0] rf_filter_coeff389_a;
	wire [7:0] rf_filter_coeff389_b;
	wire [7:0] rf_filter_coeff390_a;
	wire [7:0] rf_filter_coeff390_b;
	wire [7:0] rf_filter_coeff391_a;
	wire [7:0] rf_filter_coeff391_b;
	wire [7:0] rf_filter_coeff392_a;
	wire [7:0] rf_filter_coeff392_b;
	wire [7:0] rf_filter_coeff393_a;
	wire [7:0] rf_filter_coeff393_b;
	wire [7:0] rf_filter_coeff394_a;
	wire [7:0] rf_filter_coeff394_b;
	wire [7:0] rf_filter_coeff395_a;
	wire [7:0] rf_filter_coeff395_b;
	wire [7:0] rf_filter_coeff396_a;
	wire [7:0] rf_filter_coeff396_b;
	wire [7:0] rf_filter_coeff397_a;
	wire [7:0] rf_filter_coeff397_b;
	wire [7:0] rf_filter_coeff398_a;
	wire [7:0] rf_filter_coeff398_b;
	wire [7:0] rf_filter_coeff399_a;
	wire [7:0] rf_filter_coeff399_b;
	wire [7:0] rf_filter_coeff400_a;
	wire [7:0] rf_filter_coeff400_b;
	wire [7:0] rf_filter_coeff401_a;
	wire [7:0] rf_filter_coeff401_b;
	wire [7:0] rf_filter_coeff402_a;
	wire [7:0] rf_filter_coeff402_b;
	wire [7:0] rf_filter_coeff403_a;
	wire [7:0] rf_filter_coeff403_b;
	wire [7:0] rf_filter_coeff404_a;
	wire [7:0] rf_filter_coeff404_b;
	wire [7:0] rf_filter_coeff405_a;
	wire [7:0] rf_filter_coeff405_b;
	wire [7:0] rf_filter_coeff406_a;
	wire [7:0] rf_filter_coeff406_b;
	wire [7:0] rf_filter_coeff407_a;
	wire [7:0] rf_filter_coeff407_b;
	wire [7:0] rf_filter_coeff408_a;
	wire [7:0] rf_filter_coeff408_b;
	wire [7:0] rf_filter_coeff409_a;
	wire [7:0] rf_filter_coeff409_b;
	wire [7:0] rf_filter_coeff410_a;
	wire [7:0] rf_filter_coeff410_b;
	wire [7:0] rf_filter_coeff411_a;
	wire [7:0] rf_filter_coeff411_b;
	wire [7:0] rf_filter_coeff412_a;
	wire [7:0] rf_filter_coeff412_b;
	wire [7:0] rf_filter_coeff413_a;
	wire [7:0] rf_filter_coeff413_b;
	wire [7:0] rf_filter_coeff414_a;
	wire [7:0] rf_filter_coeff414_b;
	wire [7:0] rf_filter_coeff415_a;
	wire [7:0] rf_filter_coeff415_b;
	wire [7:0] rf_filter_coeff416_a;
	wire [7:0] rf_filter_coeff416_b;
	wire [7:0] rf_filter_coeff417_a;
	wire [7:0] rf_filter_coeff417_b;
	wire [7:0] rf_filter_coeff418_a;
	wire [7:0] rf_filter_coeff418_b;
	wire [7:0] rf_filter_coeff419_a;
	wire [7:0] rf_filter_coeff419_b;
	wire [7:0] rf_filter_coeff420_a;
	wire [7:0] rf_filter_coeff420_b;
	wire [7:0] rf_filter_coeff421_a;
	wire [7:0] rf_filter_coeff421_b;
	wire [7:0] rf_filter_coeff422_a;
	wire [7:0] rf_filter_coeff422_b;
	wire [7:0] rf_filter_coeff423_a;
	wire [7:0] rf_filter_coeff423_b;
	wire [7:0] rf_filter_coeff424_a;
	wire [7:0] rf_filter_coeff424_b;
	wire [7:0] rf_filter_coeff425_a;
	wire [7:0] rf_filter_coeff425_b;
	wire [7:0] rf_filter_coeff426_a;
	wire [7:0] rf_filter_coeff426_b;
	wire [7:0] rf_filter_coeff427_a;
	wire [7:0] rf_filter_coeff427_b;
	wire [7:0] rf_filter_coeff428_a;
	wire [7:0] rf_filter_coeff428_b;
	wire [7:0] rf_filter_coeff429_a;
	wire [7:0] rf_filter_coeff429_b;
	wire [7:0] rf_filter_coeff430_a;
	wire [7:0] rf_filter_coeff430_b;
	wire [7:0] rf_filter_coeff431_a;
	wire [7:0] rf_filter_coeff431_b;
	wire [7:0] rf_filter_coeff432_a;
	wire [7:0] rf_filter_coeff432_b;
	wire [7:0] rf_filter_coeff433_a;
	wire [7:0] rf_filter_coeff433_b;
	wire [7:0] rf_filter_coeff434_a;
	wire [7:0] rf_filter_coeff434_b;
	wire [7:0] rf_filter_coeff435_a;
	wire [7:0] rf_filter_coeff435_b;
	wire [7:0] rf_filter_coeff436_a;
	wire [7:0] rf_filter_coeff436_b;
	wire [7:0] rf_filter_coeff437_a;
	wire [7:0] rf_filter_coeff437_b;
	wire [7:0] rf_filter_coeff438_a;
	wire [7:0] rf_filter_coeff438_b;
	wire [7:0] rf_filter_coeff439_a;
	wire [7:0] rf_filter_coeff439_b;
	wire [7:0] rf_filter_coeff440_a;
	wire [7:0] rf_filter_coeff440_b;
	wire [7:0] rf_filter_coeff441_a;
	wire [7:0] rf_filter_coeff441_b;
	wire [7:0] rf_filter_coeff442_a;
	wire [7:0] rf_filter_coeff442_b;
	wire [7:0] rf_filter_coeff443_a;
	wire [7:0] rf_filter_coeff443_b;
	wire [7:0] rf_filter_coeff444_a;
	wire [7:0] rf_filter_coeff444_b;
	wire [7:0] rf_filter_coeff445_a;
	wire [7:0] rf_filter_coeff445_b;
	wire [7:0] rf_filter_coeff446_a;
	wire [7:0] rf_filter_coeff446_b;
	wire [7:0] rf_filter_coeff447_a;
	wire [7:0] rf_filter_coeff447_b;
	wire [7:0] rf_filter_coeff448_a;
	wire [7:0] rf_filter_coeff448_b;
	wire [7:0] rf_filter_coeff449_a;
	wire [7:0] rf_filter_coeff449_b;
	wire [7:0] rf_filter_coeff450_a;
	wire [7:0] rf_filter_coeff450_b;
	wire [7:0] rf_filter_coeff451_a;
	wire [7:0] rf_filter_coeff451_b;
	wire [7:0] rf_filter_coeff452_a;
	wire [7:0] rf_filter_coeff452_b;
	wire [7:0] rf_filter_coeff453_a;
	wire [7:0] rf_filter_coeff453_b;
	wire [7:0] rf_filter_coeff454_a;
	wire [7:0] rf_filter_coeff454_b;
	wire [7:0] rf_filter_coeff455_a;
	wire [7:0] rf_filter_coeff455_b;
	wire [7:0] rf_filter_coeff456_a;
	wire [7:0] rf_filter_coeff456_b;
	wire [7:0] rf_filter_coeff457_a;
	wire [7:0] rf_filter_coeff457_b;
	wire [7:0] rf_filter_coeff458_a;
	wire [7:0] rf_filter_coeff458_b;
	wire [7:0] rf_filter_coeff459_a;
	wire [7:0] rf_filter_coeff459_b;
	wire [7:0] rf_filter_coeff460_a;
	wire [7:0] rf_filter_coeff460_b;
	wire [7:0] rf_filter_coeff461_a;
	wire [7:0] rf_filter_coeff461_b;
	wire [7:0] rf_filter_coeff462_a;
	wire [7:0] rf_filter_coeff462_b;
	wire [7:0] rf_filter_coeff463_a;
	wire [7:0] rf_filter_coeff463_b;
	wire [7:0] rf_filter_coeff464_a;
	wire [7:0] rf_filter_coeff464_b;
	wire [7:0] rf_filter_coeff465_a;
	wire [7:0] rf_filter_coeff465_b;
	wire [7:0] rf_filter_coeff466_a;
	wire [7:0] rf_filter_coeff466_b;
	wire [7:0] rf_filter_coeff467_a;
	wire [7:0] rf_filter_coeff467_b;
	wire [7:0] rf_filter_coeff468_a;
	wire [7:0] rf_filter_coeff468_b;
	wire [7:0] rf_filter_coeff469_a;
	wire [7:0] rf_filter_coeff469_b;
	wire [7:0] rf_filter_coeff470_a;
	wire [7:0] rf_filter_coeff470_b;
	wire [7:0] rf_filter_coeff471_a;
	wire [7:0] rf_filter_coeff471_b;
	wire [7:0] rf_filter_coeff472_a;
	wire [7:0] rf_filter_coeff472_b;
	wire [7:0] rf_filter_coeff473_a;
	wire [7:0] rf_filter_coeff473_b;
	wire [7:0] rf_filter_coeff474_a;
	wire [7:0] rf_filter_coeff474_b;
	wire [7:0] rf_filter_coeff475_a;
	wire [7:0] rf_filter_coeff475_b;
	wire [7:0] rf_filter_coeff476_a;
	wire [7:0] rf_filter_coeff476_b;
	wire [7:0] rf_filter_coeff477_a;
	wire [7:0] rf_filter_coeff477_b;
	wire [7:0] rf_filter_coeff478_a;
	wire [7:0] rf_filter_coeff478_b;
	wire [7:0] rf_filter_coeff479_a;
	wire [7:0] rf_filter_coeff479_b;
	wire [7:0] rf_filter_coeff480_a;
	wire [7:0] rf_filter_coeff480_b;
	wire [7:0] rf_filter_coeff481_a;
	wire [7:0] rf_filter_coeff481_b;
	wire [7:0] rf_filter_coeff482_a;
	wire [7:0] rf_filter_coeff482_b;
	wire [7:0] rf_filter_coeff483_a;
	wire [7:0] rf_filter_coeff483_b;
	wire [7:0] rf_filter_coeff484_a;
	wire [7:0] rf_filter_coeff484_b;
	wire [7:0] rf_filter_coeff485_a;
	wire [7:0] rf_filter_coeff485_b;
	wire [7:0] rf_filter_coeff486_a;
	wire [7:0] rf_filter_coeff486_b;
	wire [7:0] rf_filter_coeff487_a;
	wire [7:0] rf_filter_coeff487_b;
	wire [7:0] rf_filter_coeff488_a;
	wire [7:0] rf_filter_coeff488_b;
	wire [7:0] rf_filter_coeff489_a;
	wire [7:0] rf_filter_coeff489_b;
	wire [7:0] rf_filter_coeff490_a;
	wire [7:0] rf_filter_coeff490_b;
	wire [7:0] rf_filter_coeff491_a;
	wire [7:0] rf_filter_coeff491_b;
	wire [7:0] rf_filter_coeff492_a;
	wire [7:0] rf_filter_coeff492_b;
	wire [7:0] rf_filter_coeff493_a;
	wire [7:0] rf_filter_coeff493_b;
	wire [7:0] rf_filter_coeff494_a;
	wire [7:0] rf_filter_coeff494_b;
	wire [7:0] rf_filter_coeff495_a;
	wire [7:0] rf_filter_coeff495_b;
	wire [7:0] rf_filter_coeff496_a;
	wire [7:0] rf_filter_coeff496_b;
	wire [7:0] rf_filter_coeff497_a;
	wire [7:0] rf_filter_coeff497_b;
	wire [7:0] rf_filter_coeff498_a;
	wire [7:0] rf_filter_coeff498_b;
	wire [7:0] rf_filter_coeff499_a;
	wire [7:0] rf_filter_coeff499_b;
	wire [7:0] rf_filter_coeff500_a;
	wire [7:0] rf_filter_coeff500_b;
	wire [7:0] rf_filter_coeff501_a;
	wire [7:0] rf_filter_coeff501_b;
	wire [7:0] rf_filter_coeff502_a;
	wire [7:0] rf_filter_coeff502_b;
	wire [7:0] rf_filter_coeff503_a;
	wire [7:0] rf_filter_coeff503_b;
	wire [7:0] rf_filter_coeff504_a;
	wire [7:0] rf_filter_coeff504_b;
	wire [7:0] rf_filter_coeff505_a;
	wire [7:0] rf_filter_coeff505_b;
	wire [7:0] rf_filter_coeff506_a;
	wire [7:0] rf_filter_coeff506_b;
	wire [7:0] rf_filter_coeff507_a;
	wire [7:0] rf_filter_coeff507_b;
	wire [7:0] rf_filter_coeff508_a;
	wire [7:0] rf_filter_coeff508_b;
	wire [7:0] rf_filter_coeff509_a;
	wire [7:0] rf_filter_coeff509_b;
	wire [7:0] rf_filter_coeff510_a;
	wire [7:0] rf_filter_coeff510_b;
	wire [7:0] rf_filter_coeff511_a;
	wire [7:0] rf_filter_coeff511_b;

	// Instantiate the Unit Under Test (UUT)
	register uut (
		.rst_n(rst_n), 
		.clk(clk), 
		.addr(addr), 
		.wdata(wdata), 
		.w_enable(w_enable), 
		.wxfc(wxfc), 
		.rxfc(rxfc), 
		.ro_fifo_underrun(ro_fifo_underrun), 
		.ro_fifo_overrun(ro_fifo_overrun), 
		.rdata(rdata), 
		.rf_i2si_bist_en(rf_i2si_bist_en), 
		.rf_filter_shift(rf_filter_shift), 
		.rf_filter_clip_en(rf_filter_clip_en), 
		.ro_filter_ovf_flag(ro_filter_ovf_flag), 
		.trig_fifo_overrun(trig_fifo_overrun), 
		.trig_fifo_underrun(trig_fifo_underrun), 
		.trig_filter_ovf_flag_clear(trig_filter_ovf_flag_clear), 
		.rf_i2si_bist_start_val_a(rf_i2si_bist_start_val_a), 
		.rf_i2si_bist_start_val_b(rf_i2si_bist_start_val_b), 
		.rf_i2si_bist_incr(rf_i2si_bist_incr), 
		.rf_i2si_bist_upper_limit_a(rf_i2si_bist_upper_limit_a), 
		.rf_i2si_bist_upper_limit_b(rf_i2si_bist_upper_limit_b), 
		.rf_filter_coeff0_a(rf_filter_coeff0_a), 
		.rf_filter_coeff0_b(rf_filter_coeff0_b), 
		.rf_filter_coeff1_a(rf_filter_coeff1_a), 
		.rf_filter_coeff1_b(rf_filter_coeff1_b), 
		.rf_filter_coeff2_a(rf_filter_coeff2_a), 
		.rf_filter_coeff2_b(rf_filter_coeff2_b), 
		.rf_filter_coeff3_a(rf_filter_coeff3_a), 
		.rf_filter_coeff3_b(rf_filter_coeff3_b), 
		.rf_filter_coeff4_a(rf_filter_coeff4_a), 
		.rf_filter_coeff4_b(rf_filter_coeff4_b), 
		.rf_filter_coeff5_a(rf_filter_coeff5_a), 
		.rf_filter_coeff5_b(rf_filter_coeff5_b), 
		.rf_filter_coeff6_a(rf_filter_coeff6_a), 
		.rf_filter_coeff6_b(rf_filter_coeff6_b), 
		.rf_filter_coeff7_a(rf_filter_coeff7_a), 
		.rf_filter_coeff7_b(rf_filter_coeff7_b), 
		.rf_filter_coeff8_a(rf_filter_coeff8_a), 
		.rf_filter_coeff8_b(rf_filter_coeff8_b), 
		.rf_filter_coeff9_a(rf_filter_coeff9_a), 
		.rf_filter_coeff9_b(rf_filter_coeff9_b), 
		.rf_filter_coeff10_a(rf_filter_coeff10_a), 
		.rf_filter_coeff10_b(rf_filter_coeff10_b), 
		.rf_filter_coeff11_a(rf_filter_coeff11_a), 
		.rf_filter_coeff11_b(rf_filter_coeff11_b), 
		.rf_filter_coeff12_a(rf_filter_coeff12_a), 
		.rf_filter_coeff12_b(rf_filter_coeff12_b), 
		.rf_filter_coeff13_a(rf_filter_coeff13_a), 
		.rf_filter_coeff13_b(rf_filter_coeff13_b), 
		.rf_filter_coeff14_a(rf_filter_coeff14_a), 
		.rf_filter_coeff14_b(rf_filter_coeff14_b), 
		.rf_filter_coeff15_a(rf_filter_coeff15_a), 
		.rf_filter_coeff15_b(rf_filter_coeff15_b), 
		.rf_filter_coeff16_a(rf_filter_coeff16_a), 
		.rf_filter_coeff16_b(rf_filter_coeff16_b), 
		.rf_filter_coeff17_a(rf_filter_coeff17_a), 
		.rf_filter_coeff17_b(rf_filter_coeff17_b), 
		.rf_filter_coeff18_a(rf_filter_coeff18_a), 
		.rf_filter_coeff18_b(rf_filter_coeff18_b), 
		.rf_filter_coeff19_a(rf_filter_coeff19_a), 
		.rf_filter_coeff19_b(rf_filter_coeff19_b), 
		.rf_filter_coeff20_a(rf_filter_coeff20_a), 
		.rf_filter_coeff20_b(rf_filter_coeff20_b), 
		.rf_filter_coeff21_a(rf_filter_coeff21_a), 
		.rf_filter_coeff21_b(rf_filter_coeff21_b), 
		.rf_filter_coeff22_a(rf_filter_coeff22_a), 
		.rf_filter_coeff22_b(rf_filter_coeff22_b), 
		.rf_filter_coeff23_a(rf_filter_coeff23_a), 
		.rf_filter_coeff23_b(rf_filter_coeff23_b), 
		.rf_filter_coeff24_a(rf_filter_coeff24_a), 
		.rf_filter_coeff24_b(rf_filter_coeff24_b), 
		.rf_filter_coeff25_a(rf_filter_coeff25_a), 
		.rf_filter_coeff25_b(rf_filter_coeff25_b), 
		.rf_filter_coeff26_a(rf_filter_coeff26_a), 
		.rf_filter_coeff26_b(rf_filter_coeff26_b), 
		.rf_filter_coeff27_a(rf_filter_coeff27_a), 
		.rf_filter_coeff27_b(rf_filter_coeff27_b), 
		.rf_filter_coeff28_a(rf_filter_coeff28_a), 
		.rf_filter_coeff28_b(rf_filter_coeff28_b), 
		.rf_filter_coeff29_a(rf_filter_coeff29_a), 
		.rf_filter_coeff29_b(rf_filter_coeff29_b), 
		.rf_filter_coeff30_a(rf_filter_coeff30_a), 
		.rf_filter_coeff30_b(rf_filter_coeff30_b), 
		.rf_filter_coeff31_a(rf_filter_coeff31_a), 
		.rf_filter_coeff31_b(rf_filter_coeff31_b), 
		.rf_filter_coeff32_a(rf_filter_coeff32_a), 
		.rf_filter_coeff32_b(rf_filter_coeff32_b), 
		.rf_filter_coeff33_a(rf_filter_coeff33_a), 
		.rf_filter_coeff33_b(rf_filter_coeff33_b), 
		.rf_filter_coeff34_a(rf_filter_coeff34_a), 
		.rf_filter_coeff34_b(rf_filter_coeff34_b), 
		.rf_filter_coeff35_a(rf_filter_coeff35_a), 
		.rf_filter_coeff35_b(rf_filter_coeff35_b), 
		.rf_filter_coeff36_a(rf_filter_coeff36_a), 
		.rf_filter_coeff36_b(rf_filter_coeff36_b), 
		.rf_filter_coeff37_a(rf_filter_coeff37_a), 
		.rf_filter_coeff37_b(rf_filter_coeff37_b), 
		.rf_filter_coeff38_a(rf_filter_coeff38_a), 
		.rf_filter_coeff38_b(rf_filter_coeff38_b), 
		.rf_filter_coeff39_a(rf_filter_coeff39_a), 
		.rf_filter_coeff39_b(rf_filter_coeff39_b), 
		.rf_filter_coeff40_a(rf_filter_coeff40_a), 
		.rf_filter_coeff40_b(rf_filter_coeff40_b), 
		.rf_filter_coeff41_a(rf_filter_coeff41_a), 
		.rf_filter_coeff41_b(rf_filter_coeff41_b), 
		.rf_filter_coeff42_a(rf_filter_coeff42_a), 
		.rf_filter_coeff42_b(rf_filter_coeff42_b), 
		.rf_filter_coeff43_a(rf_filter_coeff43_a), 
		.rf_filter_coeff43_b(rf_filter_coeff43_b), 
		.rf_filter_coeff44_a(rf_filter_coeff44_a), 
		.rf_filter_coeff44_b(rf_filter_coeff44_b), 
		.rf_filter_coeff45_a(rf_filter_coeff45_a), 
		.rf_filter_coeff45_b(rf_filter_coeff45_b), 
		.rf_filter_coeff46_a(rf_filter_coeff46_a), 
		.rf_filter_coeff46_b(rf_filter_coeff46_b), 
		.rf_filter_coeff47_a(rf_filter_coeff47_a), 
		.rf_filter_coeff47_b(rf_filter_coeff47_b), 
		.rf_filter_coeff48_a(rf_filter_coeff48_a), 
		.rf_filter_coeff48_b(rf_filter_coeff48_b), 
		.rf_filter_coeff49_a(rf_filter_coeff49_a), 
		.rf_filter_coeff49_b(rf_filter_coeff49_b), 
		.rf_filter_coeff50_a(rf_filter_coeff50_a), 
		.rf_filter_coeff50_b(rf_filter_coeff50_b), 
		.rf_filter_coeff51_a(rf_filter_coeff51_a), 
		.rf_filter_coeff51_b(rf_filter_coeff51_b), 
		.rf_filter_coeff52_a(rf_filter_coeff52_a), 
		.rf_filter_coeff52_b(rf_filter_coeff52_b), 
		.rf_filter_coeff53_a(rf_filter_coeff53_a), 
		.rf_filter_coeff53_b(rf_filter_coeff53_b), 
		.rf_filter_coeff54_a(rf_filter_coeff54_a), 
		.rf_filter_coeff54_b(rf_filter_coeff54_b), 
		.rf_filter_coeff55_a(rf_filter_coeff55_a), 
		.rf_filter_coeff55_b(rf_filter_coeff55_b), 
		.rf_filter_coeff56_a(rf_filter_coeff56_a), 
		.rf_filter_coeff56_b(rf_filter_coeff56_b), 
		.rf_filter_coeff57_a(rf_filter_coeff57_a), 
		.rf_filter_coeff57_b(rf_filter_coeff57_b), 
		.rf_filter_coeff58_a(rf_filter_coeff58_a), 
		.rf_filter_coeff58_b(rf_filter_coeff58_b), 
		.rf_filter_coeff59_a(rf_filter_coeff59_a), 
		.rf_filter_coeff59_b(rf_filter_coeff59_b), 
		.rf_filter_coeff60_a(rf_filter_coeff60_a), 
		.rf_filter_coeff60_b(rf_filter_coeff60_b), 
		.rf_filter_coeff61_a(rf_filter_coeff61_a), 
		.rf_filter_coeff61_b(rf_filter_coeff61_b), 
		.rf_filter_coeff62_a(rf_filter_coeff62_a), 
		.rf_filter_coeff62_b(rf_filter_coeff62_b), 
		.rf_filter_coeff63_a(rf_filter_coeff63_a), 
		.rf_filter_coeff63_b(rf_filter_coeff63_b), 
		.rf_filter_coeff64_a(rf_filter_coeff64_a), 
		.rf_filter_coeff64_b(rf_filter_coeff64_b), 
		.rf_filter_coeff65_a(rf_filter_coeff65_a), 
		.rf_filter_coeff65_b(rf_filter_coeff65_b), 
		.rf_filter_coeff66_a(rf_filter_coeff66_a), 
		.rf_filter_coeff66_b(rf_filter_coeff66_b), 
		.rf_filter_coeff67_a(rf_filter_coeff67_a), 
		.rf_filter_coeff67_b(rf_filter_coeff67_b), 
		.rf_filter_coeff68_a(rf_filter_coeff68_a), 
		.rf_filter_coeff68_b(rf_filter_coeff68_b), 
		.rf_filter_coeff69_a(rf_filter_coeff69_a), 
		.rf_filter_coeff69_b(rf_filter_coeff69_b), 
		.rf_filter_coeff70_a(rf_filter_coeff70_a), 
		.rf_filter_coeff70_b(rf_filter_coeff70_b), 
		.rf_filter_coeff71_a(rf_filter_coeff71_a), 
		.rf_filter_coeff71_b(rf_filter_coeff71_b), 
		.rf_filter_coeff72_a(rf_filter_coeff72_a), 
		.rf_filter_coeff72_b(rf_filter_coeff72_b), 
		.rf_filter_coeff73_a(rf_filter_coeff73_a), 
		.rf_filter_coeff73_b(rf_filter_coeff73_b), 
		.rf_filter_coeff74_a(rf_filter_coeff74_a), 
		.rf_filter_coeff74_b(rf_filter_coeff74_b), 
		.rf_filter_coeff75_a(rf_filter_coeff75_a), 
		.rf_filter_coeff75_b(rf_filter_coeff75_b), 
		.rf_filter_coeff76_a(rf_filter_coeff76_a), 
		.rf_filter_coeff76_b(rf_filter_coeff76_b), 
		.rf_filter_coeff77_a(rf_filter_coeff77_a), 
		.rf_filter_coeff77_b(rf_filter_coeff77_b), 
		.rf_filter_coeff78_a(rf_filter_coeff78_a), 
		.rf_filter_coeff78_b(rf_filter_coeff78_b), 
		.rf_filter_coeff79_a(rf_filter_coeff79_a), 
		.rf_filter_coeff79_b(rf_filter_coeff79_b), 
		.rf_filter_coeff80_a(rf_filter_coeff80_a), 
		.rf_filter_coeff80_b(rf_filter_coeff80_b), 
		.rf_filter_coeff81_a(rf_filter_coeff81_a), 
		.rf_filter_coeff81_b(rf_filter_coeff81_b), 
		.rf_filter_coeff82_a(rf_filter_coeff82_a), 
		.rf_filter_coeff82_b(rf_filter_coeff82_b), 
		.rf_filter_coeff83_a(rf_filter_coeff83_a), 
		.rf_filter_coeff83_b(rf_filter_coeff83_b), 
		.rf_filter_coeff84_a(rf_filter_coeff84_a), 
		.rf_filter_coeff84_b(rf_filter_coeff84_b), 
		.rf_filter_coeff85_a(rf_filter_coeff85_a), 
		.rf_filter_coeff85_b(rf_filter_coeff85_b), 
		.rf_filter_coeff86_a(rf_filter_coeff86_a), 
		.rf_filter_coeff86_b(rf_filter_coeff86_b), 
		.rf_filter_coeff87_a(rf_filter_coeff87_a), 
		.rf_filter_coeff87_b(rf_filter_coeff87_b), 
		.rf_filter_coeff88_a(rf_filter_coeff88_a), 
		.rf_filter_coeff88_b(rf_filter_coeff88_b), 
		.rf_filter_coeff89_a(rf_filter_coeff89_a), 
		.rf_filter_coeff89_b(rf_filter_coeff89_b), 
		.rf_filter_coeff90_a(rf_filter_coeff90_a), 
		.rf_filter_coeff90_b(rf_filter_coeff90_b), 
		.rf_filter_coeff91_a(rf_filter_coeff91_a), 
		.rf_filter_coeff91_b(rf_filter_coeff91_b), 
		.rf_filter_coeff92_a(rf_filter_coeff92_a), 
		.rf_filter_coeff92_b(rf_filter_coeff92_b), 
		.rf_filter_coeff93_a(rf_filter_coeff93_a), 
		.rf_filter_coeff93_b(rf_filter_coeff93_b), 
		.rf_filter_coeff94_a(rf_filter_coeff94_a), 
		.rf_filter_coeff94_b(rf_filter_coeff94_b), 
		.rf_filter_coeff95_a(rf_filter_coeff95_a), 
		.rf_filter_coeff95_b(rf_filter_coeff95_b), 
		.rf_filter_coeff96_a(rf_filter_coeff96_a), 
		.rf_filter_coeff96_b(rf_filter_coeff96_b), 
		.rf_filter_coeff97_a(rf_filter_coeff97_a), 
		.rf_filter_coeff97_b(rf_filter_coeff97_b), 
		.rf_filter_coeff98_a(rf_filter_coeff98_a), 
		.rf_filter_coeff98_b(rf_filter_coeff98_b), 
		.rf_filter_coeff99_a(rf_filter_coeff99_a), 
		.rf_filter_coeff99_b(rf_filter_coeff99_b), 
		.rf_filter_coeff100_a(rf_filter_coeff100_a), 
		.rf_filter_coeff100_b(rf_filter_coeff100_b), 
		.rf_filter_coeff101_a(rf_filter_coeff101_a), 
		.rf_filter_coeff101_b(rf_filter_coeff101_b), 
		.rf_filter_coeff102_a(rf_filter_coeff102_a), 
		.rf_filter_coeff102_b(rf_filter_coeff102_b), 
		.rf_filter_coeff103_a(rf_filter_coeff103_a), 
		.rf_filter_coeff103_b(rf_filter_coeff103_b), 
		.rf_filter_coeff104_a(rf_filter_coeff104_a), 
		.rf_filter_coeff104_b(rf_filter_coeff104_b), 
		.rf_filter_coeff105_a(rf_filter_coeff105_a), 
		.rf_filter_coeff105_b(rf_filter_coeff105_b), 
		.rf_filter_coeff106_a(rf_filter_coeff106_a), 
		.rf_filter_coeff106_b(rf_filter_coeff106_b), 
		.rf_filter_coeff107_a(rf_filter_coeff107_a), 
		.rf_filter_coeff107_b(rf_filter_coeff107_b), 
		.rf_filter_coeff108_a(rf_filter_coeff108_a), 
		.rf_filter_coeff108_b(rf_filter_coeff108_b), 
		.rf_filter_coeff109_a(rf_filter_coeff109_a), 
		.rf_filter_coeff109_b(rf_filter_coeff109_b), 
		.rf_filter_coeff110_a(rf_filter_coeff110_a), 
		.rf_filter_coeff110_b(rf_filter_coeff110_b), 
		.rf_filter_coeff111_a(rf_filter_coeff111_a), 
		.rf_filter_coeff111_b(rf_filter_coeff111_b), 
		.rf_filter_coeff112_a(rf_filter_coeff112_a), 
		.rf_filter_coeff112_b(rf_filter_coeff112_b), 
		.rf_filter_coeff113_a(rf_filter_coeff113_a), 
		.rf_filter_coeff113_b(rf_filter_coeff113_b), 
		.rf_filter_coeff114_a(rf_filter_coeff114_a), 
		.rf_filter_coeff114_b(rf_filter_coeff114_b), 
		.rf_filter_coeff115_a(rf_filter_coeff115_a), 
		.rf_filter_coeff115_b(rf_filter_coeff115_b), 
		.rf_filter_coeff116_a(rf_filter_coeff116_a), 
		.rf_filter_coeff116_b(rf_filter_coeff116_b), 
		.rf_filter_coeff117_a(rf_filter_coeff117_a), 
		.rf_filter_coeff117_b(rf_filter_coeff117_b), 
		.rf_filter_coeff118_a(rf_filter_coeff118_a), 
		.rf_filter_coeff118_b(rf_filter_coeff118_b), 
		.rf_filter_coeff119_a(rf_filter_coeff119_a), 
		.rf_filter_coeff119_b(rf_filter_coeff119_b), 
		.rf_filter_coeff120_a(rf_filter_coeff120_a), 
		.rf_filter_coeff120_b(rf_filter_coeff120_b), 
		.rf_filter_coeff121_a(rf_filter_coeff121_a), 
		.rf_filter_coeff121_b(rf_filter_coeff121_b), 
		.rf_filter_coeff122_a(rf_filter_coeff122_a), 
		.rf_filter_coeff122_b(rf_filter_coeff122_b), 
		.rf_filter_coeff123_a(rf_filter_coeff123_a), 
		.rf_filter_coeff123_b(rf_filter_coeff123_b), 
		.rf_filter_coeff124_a(rf_filter_coeff124_a), 
		.rf_filter_coeff124_b(rf_filter_coeff124_b), 
		.rf_filter_coeff125_a(rf_filter_coeff125_a), 
		.rf_filter_coeff125_b(rf_filter_coeff125_b), 
		.rf_filter_coeff126_a(rf_filter_coeff126_a), 
		.rf_filter_coeff126_b(rf_filter_coeff126_b), 
		.rf_filter_coeff127_a(rf_filter_coeff127_a), 
		.rf_filter_coeff127_b(rf_filter_coeff127_b), 
		.rf_filter_coeff128_a(rf_filter_coeff128_a), 
		.rf_filter_coeff128_b(rf_filter_coeff128_b), 
		.rf_filter_coeff129_a(rf_filter_coeff129_a), 
		.rf_filter_coeff129_b(rf_filter_coeff129_b), 
		.rf_filter_coeff130_a(rf_filter_coeff130_a), 
		.rf_filter_coeff130_b(rf_filter_coeff130_b), 
		.rf_filter_coeff131_a(rf_filter_coeff131_a), 
		.rf_filter_coeff131_b(rf_filter_coeff131_b), 
		.rf_filter_coeff132_a(rf_filter_coeff132_a), 
		.rf_filter_coeff132_b(rf_filter_coeff132_b), 
		.rf_filter_coeff133_a(rf_filter_coeff133_a), 
		.rf_filter_coeff133_b(rf_filter_coeff133_b), 
		.rf_filter_coeff134_a(rf_filter_coeff134_a), 
		.rf_filter_coeff134_b(rf_filter_coeff134_b), 
		.rf_filter_coeff135_a(rf_filter_coeff135_a), 
		.rf_filter_coeff135_b(rf_filter_coeff135_b), 
		.rf_filter_coeff136_a(rf_filter_coeff136_a), 
		.rf_filter_coeff136_b(rf_filter_coeff136_b), 
		.rf_filter_coeff137_a(rf_filter_coeff137_a), 
		.rf_filter_coeff137_b(rf_filter_coeff137_b), 
		.rf_filter_coeff138_a(rf_filter_coeff138_a), 
		.rf_filter_coeff138_b(rf_filter_coeff138_b), 
		.rf_filter_coeff139_a(rf_filter_coeff139_a), 
		.rf_filter_coeff139_b(rf_filter_coeff139_b), 
		.rf_filter_coeff140_a(rf_filter_coeff140_a), 
		.rf_filter_coeff140_b(rf_filter_coeff140_b), 
		.rf_filter_coeff141_a(rf_filter_coeff141_a), 
		.rf_filter_coeff141_b(rf_filter_coeff141_b), 
		.rf_filter_coeff142_a(rf_filter_coeff142_a), 
		.rf_filter_coeff142_b(rf_filter_coeff142_b), 
		.rf_filter_coeff143_a(rf_filter_coeff143_a), 
		.rf_filter_coeff143_b(rf_filter_coeff143_b), 
		.rf_filter_coeff144_a(rf_filter_coeff144_a), 
		.rf_filter_coeff144_b(rf_filter_coeff144_b), 
		.rf_filter_coeff145_a(rf_filter_coeff145_a), 
		.rf_filter_coeff145_b(rf_filter_coeff145_b), 
		.rf_filter_coeff146_a(rf_filter_coeff146_a), 
		.rf_filter_coeff146_b(rf_filter_coeff146_b), 
		.rf_filter_coeff147_a(rf_filter_coeff147_a), 
		.rf_filter_coeff147_b(rf_filter_coeff147_b), 
		.rf_filter_coeff148_a(rf_filter_coeff148_a), 
		.rf_filter_coeff148_b(rf_filter_coeff148_b), 
		.rf_filter_coeff149_a(rf_filter_coeff149_a), 
		.rf_filter_coeff149_b(rf_filter_coeff149_b), 
		.rf_filter_coeff150_a(rf_filter_coeff150_a), 
		.rf_filter_coeff150_b(rf_filter_coeff150_b), 
		.rf_filter_coeff151_a(rf_filter_coeff151_a), 
		.rf_filter_coeff151_b(rf_filter_coeff151_b), 
		.rf_filter_coeff152_a(rf_filter_coeff152_a), 
		.rf_filter_coeff152_b(rf_filter_coeff152_b), 
		.rf_filter_coeff153_a(rf_filter_coeff153_a), 
		.rf_filter_coeff153_b(rf_filter_coeff153_b), 
		.rf_filter_coeff154_a(rf_filter_coeff154_a), 
		.rf_filter_coeff154_b(rf_filter_coeff154_b), 
		.rf_filter_coeff155_a(rf_filter_coeff155_a), 
		.rf_filter_coeff155_b(rf_filter_coeff155_b), 
		.rf_filter_coeff156_a(rf_filter_coeff156_a), 
		.rf_filter_coeff156_b(rf_filter_coeff156_b), 
		.rf_filter_coeff157_a(rf_filter_coeff157_a), 
		.rf_filter_coeff157_b(rf_filter_coeff157_b), 
		.rf_filter_coeff158_a(rf_filter_coeff158_a), 
		.rf_filter_coeff158_b(rf_filter_coeff158_b), 
		.rf_filter_coeff159_a(rf_filter_coeff159_a), 
		.rf_filter_coeff159_b(rf_filter_coeff159_b), 
		.rf_filter_coeff160_a(rf_filter_coeff160_a), 
		.rf_filter_coeff160_b(rf_filter_coeff160_b), 
		.rf_filter_coeff161_a(rf_filter_coeff161_a), 
		.rf_filter_coeff161_b(rf_filter_coeff161_b), 
		.rf_filter_coeff162_a(rf_filter_coeff162_a), 
		.rf_filter_coeff162_b(rf_filter_coeff162_b), 
		.rf_filter_coeff163_a(rf_filter_coeff163_a), 
		.rf_filter_coeff163_b(rf_filter_coeff163_b), 
		.rf_filter_coeff164_a(rf_filter_coeff164_a), 
		.rf_filter_coeff164_b(rf_filter_coeff164_b), 
		.rf_filter_coeff165_a(rf_filter_coeff165_a), 
		.rf_filter_coeff165_b(rf_filter_coeff165_b), 
		.rf_filter_coeff166_a(rf_filter_coeff166_a), 
		.rf_filter_coeff166_b(rf_filter_coeff166_b), 
		.rf_filter_coeff167_a(rf_filter_coeff167_a), 
		.rf_filter_coeff167_b(rf_filter_coeff167_b), 
		.rf_filter_coeff168_a(rf_filter_coeff168_a), 
		.rf_filter_coeff168_b(rf_filter_coeff168_b), 
		.rf_filter_coeff169_a(rf_filter_coeff169_a), 
		.rf_filter_coeff169_b(rf_filter_coeff169_b), 
		.rf_filter_coeff170_a(rf_filter_coeff170_a), 
		.rf_filter_coeff170_b(rf_filter_coeff170_b), 
		.rf_filter_coeff171_a(rf_filter_coeff171_a), 
		.rf_filter_coeff171_b(rf_filter_coeff171_b), 
		.rf_filter_coeff172_a(rf_filter_coeff172_a), 
		.rf_filter_coeff172_b(rf_filter_coeff172_b), 
		.rf_filter_coeff173_a(rf_filter_coeff173_a), 
		.rf_filter_coeff173_b(rf_filter_coeff173_b), 
		.rf_filter_coeff174_a(rf_filter_coeff174_a), 
		.rf_filter_coeff174_b(rf_filter_coeff174_b), 
		.rf_filter_coeff175_a(rf_filter_coeff175_a), 
		.rf_filter_coeff175_b(rf_filter_coeff175_b), 
		.rf_filter_coeff176_a(rf_filter_coeff176_a), 
		.rf_filter_coeff176_b(rf_filter_coeff176_b), 
		.rf_filter_coeff177_a(rf_filter_coeff177_a), 
		.rf_filter_coeff177_b(rf_filter_coeff177_b), 
		.rf_filter_coeff178_a(rf_filter_coeff178_a), 
		.rf_filter_coeff178_b(rf_filter_coeff178_b), 
		.rf_filter_coeff179_a(rf_filter_coeff179_a), 
		.rf_filter_coeff179_b(rf_filter_coeff179_b), 
		.rf_filter_coeff180_a(rf_filter_coeff180_a), 
		.rf_filter_coeff180_b(rf_filter_coeff180_b), 
		.rf_filter_coeff181_a(rf_filter_coeff181_a), 
		.rf_filter_coeff181_b(rf_filter_coeff181_b), 
		.rf_filter_coeff182_a(rf_filter_coeff182_a), 
		.rf_filter_coeff182_b(rf_filter_coeff182_b), 
		.rf_filter_coeff183_a(rf_filter_coeff183_a), 
		.rf_filter_coeff183_b(rf_filter_coeff183_b), 
		.rf_filter_coeff184_a(rf_filter_coeff184_a), 
		.rf_filter_coeff184_b(rf_filter_coeff184_b), 
		.rf_filter_coeff185_a(rf_filter_coeff185_a), 
		.rf_filter_coeff185_b(rf_filter_coeff185_b), 
		.rf_filter_coeff186_a(rf_filter_coeff186_a), 
		.rf_filter_coeff186_b(rf_filter_coeff186_b), 
		.rf_filter_coeff187_a(rf_filter_coeff187_a), 
		.rf_filter_coeff187_b(rf_filter_coeff187_b), 
		.rf_filter_coeff188_a(rf_filter_coeff188_a), 
		.rf_filter_coeff188_b(rf_filter_coeff188_b), 
		.rf_filter_coeff189_a(rf_filter_coeff189_a), 
		.rf_filter_coeff189_b(rf_filter_coeff189_b), 
		.rf_filter_coeff190_a(rf_filter_coeff190_a), 
		.rf_filter_coeff190_b(rf_filter_coeff190_b), 
		.rf_filter_coeff191_a(rf_filter_coeff191_a), 
		.rf_filter_coeff191_b(rf_filter_coeff191_b), 
		.rf_filter_coeff192_a(rf_filter_coeff192_a), 
		.rf_filter_coeff192_b(rf_filter_coeff192_b), 
		.rf_filter_coeff193_a(rf_filter_coeff193_a), 
		.rf_filter_coeff193_b(rf_filter_coeff193_b), 
		.rf_filter_coeff194_a(rf_filter_coeff194_a), 
		.rf_filter_coeff194_b(rf_filter_coeff194_b), 
		.rf_filter_coeff195_a(rf_filter_coeff195_a), 
		.rf_filter_coeff195_b(rf_filter_coeff195_b), 
		.rf_filter_coeff196_a(rf_filter_coeff196_a), 
		.rf_filter_coeff196_b(rf_filter_coeff196_b), 
		.rf_filter_coeff197_a(rf_filter_coeff197_a), 
		.rf_filter_coeff197_b(rf_filter_coeff197_b), 
		.rf_filter_coeff198_a(rf_filter_coeff198_a), 
		.rf_filter_coeff198_b(rf_filter_coeff198_b), 
		.rf_filter_coeff199_a(rf_filter_coeff199_a), 
		.rf_filter_coeff199_b(rf_filter_coeff199_b), 
		.rf_filter_coeff200_a(rf_filter_coeff200_a), 
		.rf_filter_coeff200_b(rf_filter_coeff200_b), 
		.rf_filter_coeff201_a(rf_filter_coeff201_a), 
		.rf_filter_coeff201_b(rf_filter_coeff201_b), 
		.rf_filter_coeff202_a(rf_filter_coeff202_a), 
		.rf_filter_coeff202_b(rf_filter_coeff202_b), 
		.rf_filter_coeff203_a(rf_filter_coeff203_a), 
		.rf_filter_coeff203_b(rf_filter_coeff203_b), 
		.rf_filter_coeff204_a(rf_filter_coeff204_a), 
		.rf_filter_coeff204_b(rf_filter_coeff204_b), 
		.rf_filter_coeff205_a(rf_filter_coeff205_a), 
		.rf_filter_coeff205_b(rf_filter_coeff205_b), 
		.rf_filter_coeff206_a(rf_filter_coeff206_a), 
		.rf_filter_coeff206_b(rf_filter_coeff206_b), 
		.rf_filter_coeff207_a(rf_filter_coeff207_a), 
		.rf_filter_coeff207_b(rf_filter_coeff207_b), 
		.rf_filter_coeff208_a(rf_filter_coeff208_a), 
		.rf_filter_coeff208_b(rf_filter_coeff208_b), 
		.rf_filter_coeff209_a(rf_filter_coeff209_a), 
		.rf_filter_coeff209_b(rf_filter_coeff209_b), 
		.rf_filter_coeff210_a(rf_filter_coeff210_a), 
		.rf_filter_coeff210_b(rf_filter_coeff210_b), 
		.rf_filter_coeff211_a(rf_filter_coeff211_a), 
		.rf_filter_coeff211_b(rf_filter_coeff211_b), 
		.rf_filter_coeff212_a(rf_filter_coeff212_a), 
		.rf_filter_coeff212_b(rf_filter_coeff212_b), 
		.rf_filter_coeff213_a(rf_filter_coeff213_a), 
		.rf_filter_coeff213_b(rf_filter_coeff213_b), 
		.rf_filter_coeff214_a(rf_filter_coeff214_a), 
		.rf_filter_coeff214_b(rf_filter_coeff214_b), 
		.rf_filter_coeff215_a(rf_filter_coeff215_a), 
		.rf_filter_coeff215_b(rf_filter_coeff215_b), 
		.rf_filter_coeff216_a(rf_filter_coeff216_a), 
		.rf_filter_coeff216_b(rf_filter_coeff216_b), 
		.rf_filter_coeff217_a(rf_filter_coeff217_a), 
		.rf_filter_coeff217_b(rf_filter_coeff217_b), 
		.rf_filter_coeff218_a(rf_filter_coeff218_a), 
		.rf_filter_coeff218_b(rf_filter_coeff218_b), 
		.rf_filter_coeff219_a(rf_filter_coeff219_a), 
		.rf_filter_coeff219_b(rf_filter_coeff219_b), 
		.rf_filter_coeff220_a(rf_filter_coeff220_a), 
		.rf_filter_coeff220_b(rf_filter_coeff220_b), 
		.rf_filter_coeff221_a(rf_filter_coeff221_a), 
		.rf_filter_coeff221_b(rf_filter_coeff221_b), 
		.rf_filter_coeff222_a(rf_filter_coeff222_a), 
		.rf_filter_coeff222_b(rf_filter_coeff222_b), 
		.rf_filter_coeff223_a(rf_filter_coeff223_a), 
		.rf_filter_coeff223_b(rf_filter_coeff223_b), 
		.rf_filter_coeff224_a(rf_filter_coeff224_a), 
		.rf_filter_coeff224_b(rf_filter_coeff224_b), 
		.rf_filter_coeff225_a(rf_filter_coeff225_a), 
		.rf_filter_coeff225_b(rf_filter_coeff225_b), 
		.rf_filter_coeff226_a(rf_filter_coeff226_a), 
		.rf_filter_coeff226_b(rf_filter_coeff226_b), 
		.rf_filter_coeff227_a(rf_filter_coeff227_a), 
		.rf_filter_coeff227_b(rf_filter_coeff227_b), 
		.rf_filter_coeff228_a(rf_filter_coeff228_a), 
		.rf_filter_coeff228_b(rf_filter_coeff228_b), 
		.rf_filter_coeff229_a(rf_filter_coeff229_a), 
		.rf_filter_coeff229_b(rf_filter_coeff229_b), 
		.rf_filter_coeff230_a(rf_filter_coeff230_a), 
		.rf_filter_coeff230_b(rf_filter_coeff230_b), 
		.rf_filter_coeff231_a(rf_filter_coeff231_a), 
		.rf_filter_coeff231_b(rf_filter_coeff231_b), 
		.rf_filter_coeff232_a(rf_filter_coeff232_a), 
		.rf_filter_coeff232_b(rf_filter_coeff232_b), 
		.rf_filter_coeff233_a(rf_filter_coeff233_a), 
		.rf_filter_coeff233_b(rf_filter_coeff233_b), 
		.rf_filter_coeff234_a(rf_filter_coeff234_a), 
		.rf_filter_coeff234_b(rf_filter_coeff234_b), 
		.rf_filter_coeff235_a(rf_filter_coeff235_a), 
		.rf_filter_coeff235_b(rf_filter_coeff235_b), 
		.rf_filter_coeff236_a(rf_filter_coeff236_a), 
		.rf_filter_coeff236_b(rf_filter_coeff236_b), 
		.rf_filter_coeff237_a(rf_filter_coeff237_a), 
		.rf_filter_coeff237_b(rf_filter_coeff237_b), 
		.rf_filter_coeff238_a(rf_filter_coeff238_a), 
		.rf_filter_coeff238_b(rf_filter_coeff238_b), 
		.rf_filter_coeff239_a(rf_filter_coeff239_a), 
		.rf_filter_coeff239_b(rf_filter_coeff239_b), 
		.rf_filter_coeff240_a(rf_filter_coeff240_a), 
		.rf_filter_coeff240_b(rf_filter_coeff240_b), 
		.rf_filter_coeff241_a(rf_filter_coeff241_a), 
		.rf_filter_coeff241_b(rf_filter_coeff241_b), 
		.rf_filter_coeff242_a(rf_filter_coeff242_a), 
		.rf_filter_coeff242_b(rf_filter_coeff242_b), 
		.rf_filter_coeff243_a(rf_filter_coeff243_a), 
		.rf_filter_coeff243_b(rf_filter_coeff243_b), 
		.rf_filter_coeff244_a(rf_filter_coeff244_a), 
		.rf_filter_coeff244_b(rf_filter_coeff244_b), 
		.rf_filter_coeff245_a(rf_filter_coeff245_a), 
		.rf_filter_coeff245_b(rf_filter_coeff245_b), 
		.rf_filter_coeff246_a(rf_filter_coeff246_a), 
		.rf_filter_coeff246_b(rf_filter_coeff246_b), 
		.rf_filter_coeff247_a(rf_filter_coeff247_a), 
		.rf_filter_coeff247_b(rf_filter_coeff247_b), 
		.rf_filter_coeff248_a(rf_filter_coeff248_a), 
		.rf_filter_coeff248_b(rf_filter_coeff248_b), 
		.rf_filter_coeff249_a(rf_filter_coeff249_a), 
		.rf_filter_coeff249_b(rf_filter_coeff249_b), 
		.rf_filter_coeff250_a(rf_filter_coeff250_a), 
		.rf_filter_coeff250_b(rf_filter_coeff250_b), 
		.rf_filter_coeff251_a(rf_filter_coeff251_a), 
		.rf_filter_coeff251_b(rf_filter_coeff251_b), 
		.rf_filter_coeff252_a(rf_filter_coeff252_a), 
		.rf_filter_coeff252_b(rf_filter_coeff252_b), 
		.rf_filter_coeff253_a(rf_filter_coeff253_a), 
		.rf_filter_coeff253_b(rf_filter_coeff253_b), 
		.rf_filter_coeff254_a(rf_filter_coeff254_a), 
		.rf_filter_coeff254_b(rf_filter_coeff254_b), 
		.rf_filter_coeff255_a(rf_filter_coeff255_a), 
		.rf_filter_coeff255_b(rf_filter_coeff255_b), 
		.rf_filter_coeff256_a(rf_filter_coeff256_a), 
		.rf_filter_coeff256_b(rf_filter_coeff256_b), 
		.rf_filter_coeff257_a(rf_filter_coeff257_a), 
		.rf_filter_coeff257_b(rf_filter_coeff257_b), 
		.rf_filter_coeff258_a(rf_filter_coeff258_a), 
		.rf_filter_coeff258_b(rf_filter_coeff258_b), 
		.rf_filter_coeff259_a(rf_filter_coeff259_a), 
		.rf_filter_coeff259_b(rf_filter_coeff259_b), 
		.rf_filter_coeff260_a(rf_filter_coeff260_a), 
		.rf_filter_coeff260_b(rf_filter_coeff260_b), 
		.rf_filter_coeff261_a(rf_filter_coeff261_a), 
		.rf_filter_coeff261_b(rf_filter_coeff261_b), 
		.rf_filter_coeff262_a(rf_filter_coeff262_a), 
		.rf_filter_coeff262_b(rf_filter_coeff262_b), 
		.rf_filter_coeff263_a(rf_filter_coeff263_a), 
		.rf_filter_coeff263_b(rf_filter_coeff263_b), 
		.rf_filter_coeff264_a(rf_filter_coeff264_a), 
		.rf_filter_coeff264_b(rf_filter_coeff264_b), 
		.rf_filter_coeff265_a(rf_filter_coeff265_a), 
		.rf_filter_coeff265_b(rf_filter_coeff265_b), 
		.rf_filter_coeff266_a(rf_filter_coeff266_a), 
		.rf_filter_coeff266_b(rf_filter_coeff266_b), 
		.rf_filter_coeff267_a(rf_filter_coeff267_a), 
		.rf_filter_coeff267_b(rf_filter_coeff267_b), 
		.rf_filter_coeff268_a(rf_filter_coeff268_a), 
		.rf_filter_coeff268_b(rf_filter_coeff268_b), 
		.rf_filter_coeff269_a(rf_filter_coeff269_a), 
		.rf_filter_coeff269_b(rf_filter_coeff269_b), 
		.rf_filter_coeff270_a(rf_filter_coeff270_a), 
		.rf_filter_coeff270_b(rf_filter_coeff270_b), 
		.rf_filter_coeff271_a(rf_filter_coeff271_a), 
		.rf_filter_coeff271_b(rf_filter_coeff271_b), 
		.rf_filter_coeff272_a(rf_filter_coeff272_a), 
		.rf_filter_coeff272_b(rf_filter_coeff272_b), 
		.rf_filter_coeff273_a(rf_filter_coeff273_a), 
		.rf_filter_coeff273_b(rf_filter_coeff273_b), 
		.rf_filter_coeff274_a(rf_filter_coeff274_a), 
		.rf_filter_coeff274_b(rf_filter_coeff274_b), 
		.rf_filter_coeff275_a(rf_filter_coeff275_a), 
		.rf_filter_coeff275_b(rf_filter_coeff275_b), 
		.rf_filter_coeff276_a(rf_filter_coeff276_a), 
		.rf_filter_coeff276_b(rf_filter_coeff276_b), 
		.rf_filter_coeff277_a(rf_filter_coeff277_a), 
		.rf_filter_coeff277_b(rf_filter_coeff277_b), 
		.rf_filter_coeff278_a(rf_filter_coeff278_a), 
		.rf_filter_coeff278_b(rf_filter_coeff278_b), 
		.rf_filter_coeff279_a(rf_filter_coeff279_a), 
		.rf_filter_coeff279_b(rf_filter_coeff279_b), 
		.rf_filter_coeff280_a(rf_filter_coeff280_a), 
		.rf_filter_coeff280_b(rf_filter_coeff280_b), 
		.rf_filter_coeff281_a(rf_filter_coeff281_a), 
		.rf_filter_coeff281_b(rf_filter_coeff281_b), 
		.rf_filter_coeff282_a(rf_filter_coeff282_a), 
		.rf_filter_coeff282_b(rf_filter_coeff282_b), 
		.rf_filter_coeff283_a(rf_filter_coeff283_a), 
		.rf_filter_coeff283_b(rf_filter_coeff283_b), 
		.rf_filter_coeff284_a(rf_filter_coeff284_a), 
		.rf_filter_coeff284_b(rf_filter_coeff284_b), 
		.rf_filter_coeff285_a(rf_filter_coeff285_a), 
		.rf_filter_coeff285_b(rf_filter_coeff285_b), 
		.rf_filter_coeff286_a(rf_filter_coeff286_a), 
		.rf_filter_coeff286_b(rf_filter_coeff286_b), 
		.rf_filter_coeff287_a(rf_filter_coeff287_a), 
		.rf_filter_coeff287_b(rf_filter_coeff287_b), 
		.rf_filter_coeff288_a(rf_filter_coeff288_a), 
		.rf_filter_coeff288_b(rf_filter_coeff288_b), 
		.rf_filter_coeff289_a(rf_filter_coeff289_a), 
		.rf_filter_coeff289_b(rf_filter_coeff289_b), 
		.rf_filter_coeff290_a(rf_filter_coeff290_a), 
		.rf_filter_coeff290_b(rf_filter_coeff290_b), 
		.rf_filter_coeff291_a(rf_filter_coeff291_a), 
		.rf_filter_coeff291_b(rf_filter_coeff291_b), 
		.rf_filter_coeff292_a(rf_filter_coeff292_a), 
		.rf_filter_coeff292_b(rf_filter_coeff292_b), 
		.rf_filter_coeff293_a(rf_filter_coeff293_a), 
		.rf_filter_coeff293_b(rf_filter_coeff293_b), 
		.rf_filter_coeff294_a(rf_filter_coeff294_a), 
		.rf_filter_coeff294_b(rf_filter_coeff294_b), 
		.rf_filter_coeff295_a(rf_filter_coeff295_a), 
		.rf_filter_coeff295_b(rf_filter_coeff295_b), 
		.rf_filter_coeff296_a(rf_filter_coeff296_a), 
		.rf_filter_coeff296_b(rf_filter_coeff296_b), 
		.rf_filter_coeff297_a(rf_filter_coeff297_a), 
		.rf_filter_coeff297_b(rf_filter_coeff297_b), 
		.rf_filter_coeff298_a(rf_filter_coeff298_a), 
		.rf_filter_coeff298_b(rf_filter_coeff298_b), 
		.rf_filter_coeff299_a(rf_filter_coeff299_a), 
		.rf_filter_coeff299_b(rf_filter_coeff299_b), 
		.rf_filter_coeff300_a(rf_filter_coeff300_a), 
		.rf_filter_coeff300_b(rf_filter_coeff300_b), 
		.rf_filter_coeff301_a(rf_filter_coeff301_a), 
		.rf_filter_coeff301_b(rf_filter_coeff301_b), 
		.rf_filter_coeff302_a(rf_filter_coeff302_a), 
		.rf_filter_coeff302_b(rf_filter_coeff302_b), 
		.rf_filter_coeff303_a(rf_filter_coeff303_a), 
		.rf_filter_coeff303_b(rf_filter_coeff303_b), 
		.rf_filter_coeff304_a(rf_filter_coeff304_a), 
		.rf_filter_coeff304_b(rf_filter_coeff304_b), 
		.rf_filter_coeff305_a(rf_filter_coeff305_a), 
		.rf_filter_coeff305_b(rf_filter_coeff305_b), 
		.rf_filter_coeff306_a(rf_filter_coeff306_a), 
		.rf_filter_coeff306_b(rf_filter_coeff306_b), 
		.rf_filter_coeff307_a(rf_filter_coeff307_a), 
		.rf_filter_coeff307_b(rf_filter_coeff307_b), 
		.rf_filter_coeff308_a(rf_filter_coeff308_a), 
		.rf_filter_coeff308_b(rf_filter_coeff308_b), 
		.rf_filter_coeff309_a(rf_filter_coeff309_a), 
		.rf_filter_coeff309_b(rf_filter_coeff309_b), 
		.rf_filter_coeff310_a(rf_filter_coeff310_a), 
		.rf_filter_coeff310_b(rf_filter_coeff310_b), 
		.rf_filter_coeff311_a(rf_filter_coeff311_a), 
		.rf_filter_coeff311_b(rf_filter_coeff311_b), 
		.rf_filter_coeff312_a(rf_filter_coeff312_a), 
		.rf_filter_coeff312_b(rf_filter_coeff312_b), 
		.rf_filter_coeff313_a(rf_filter_coeff313_a), 
		.rf_filter_coeff313_b(rf_filter_coeff313_b), 
		.rf_filter_coeff314_a(rf_filter_coeff314_a), 
		.rf_filter_coeff314_b(rf_filter_coeff314_b), 
		.rf_filter_coeff315_a(rf_filter_coeff315_a), 
		.rf_filter_coeff315_b(rf_filter_coeff315_b), 
		.rf_filter_coeff316_a(rf_filter_coeff316_a), 
		.rf_filter_coeff316_b(rf_filter_coeff316_b), 
		.rf_filter_coeff317_a(rf_filter_coeff317_a), 
		.rf_filter_coeff317_b(rf_filter_coeff317_b), 
		.rf_filter_coeff318_a(rf_filter_coeff318_a), 
		.rf_filter_coeff318_b(rf_filter_coeff318_b), 
		.rf_filter_coeff319_a(rf_filter_coeff319_a), 
		.rf_filter_coeff319_b(rf_filter_coeff319_b), 
		.rf_filter_coeff320_a(rf_filter_coeff320_a), 
		.rf_filter_coeff320_b(rf_filter_coeff320_b), 
		.rf_filter_coeff321_a(rf_filter_coeff321_a), 
		.rf_filter_coeff321_b(rf_filter_coeff321_b), 
		.rf_filter_coeff322_a(rf_filter_coeff322_a), 
		.rf_filter_coeff322_b(rf_filter_coeff322_b), 
		.rf_filter_coeff323_a(rf_filter_coeff323_a), 
		.rf_filter_coeff323_b(rf_filter_coeff323_b), 
		.rf_filter_coeff324_a(rf_filter_coeff324_a), 
		.rf_filter_coeff324_b(rf_filter_coeff324_b), 
		.rf_filter_coeff325_a(rf_filter_coeff325_a), 
		.rf_filter_coeff325_b(rf_filter_coeff325_b), 
		.rf_filter_coeff326_a(rf_filter_coeff326_a), 
		.rf_filter_coeff326_b(rf_filter_coeff326_b), 
		.rf_filter_coeff327_a(rf_filter_coeff327_a), 
		.rf_filter_coeff327_b(rf_filter_coeff327_b), 
		.rf_filter_coeff328_a(rf_filter_coeff328_a), 
		.rf_filter_coeff328_b(rf_filter_coeff328_b), 
		.rf_filter_coeff329_a(rf_filter_coeff329_a), 
		.rf_filter_coeff329_b(rf_filter_coeff329_b), 
		.rf_filter_coeff330_a(rf_filter_coeff330_a), 
		.rf_filter_coeff330_b(rf_filter_coeff330_b), 
		.rf_filter_coeff331_a(rf_filter_coeff331_a), 
		.rf_filter_coeff331_b(rf_filter_coeff331_b), 
		.rf_filter_coeff332_a(rf_filter_coeff332_a), 
		.rf_filter_coeff332_b(rf_filter_coeff332_b), 
		.rf_filter_coeff333_a(rf_filter_coeff333_a), 
		.rf_filter_coeff333_b(rf_filter_coeff333_b), 
		.rf_filter_coeff334_a(rf_filter_coeff334_a), 
		.rf_filter_coeff334_b(rf_filter_coeff334_b), 
		.rf_filter_coeff335_a(rf_filter_coeff335_a), 
		.rf_filter_coeff335_b(rf_filter_coeff335_b), 
		.rf_filter_coeff336_a(rf_filter_coeff336_a), 
		.rf_filter_coeff336_b(rf_filter_coeff336_b), 
		.rf_filter_coeff337_a(rf_filter_coeff337_a), 
		.rf_filter_coeff337_b(rf_filter_coeff337_b), 
		.rf_filter_coeff338_a(rf_filter_coeff338_a), 
		.rf_filter_coeff338_b(rf_filter_coeff338_b), 
		.rf_filter_coeff339_a(rf_filter_coeff339_a), 
		.rf_filter_coeff339_b(rf_filter_coeff339_b), 
		.rf_filter_coeff340_a(rf_filter_coeff340_a), 
		.rf_filter_coeff340_b(rf_filter_coeff340_b), 
		.rf_filter_coeff341_a(rf_filter_coeff341_a), 
		.rf_filter_coeff341_b(rf_filter_coeff341_b), 
		.rf_filter_coeff342_a(rf_filter_coeff342_a), 
		.rf_filter_coeff342_b(rf_filter_coeff342_b), 
		.rf_filter_coeff343_a(rf_filter_coeff343_a), 
		.rf_filter_coeff343_b(rf_filter_coeff343_b), 
		.rf_filter_coeff344_a(rf_filter_coeff344_a), 
		.rf_filter_coeff344_b(rf_filter_coeff344_b), 
		.rf_filter_coeff345_a(rf_filter_coeff345_a), 
		.rf_filter_coeff345_b(rf_filter_coeff345_b), 
		.rf_filter_coeff346_a(rf_filter_coeff346_a), 
		.rf_filter_coeff346_b(rf_filter_coeff346_b), 
		.rf_filter_coeff347_a(rf_filter_coeff347_a), 
		.rf_filter_coeff347_b(rf_filter_coeff347_b), 
		.rf_filter_coeff348_a(rf_filter_coeff348_a), 
		.rf_filter_coeff348_b(rf_filter_coeff348_b), 
		.rf_filter_coeff349_a(rf_filter_coeff349_a), 
		.rf_filter_coeff349_b(rf_filter_coeff349_b), 
		.rf_filter_coeff350_a(rf_filter_coeff350_a), 
		.rf_filter_coeff350_b(rf_filter_coeff350_b), 
		.rf_filter_coeff351_a(rf_filter_coeff351_a), 
		.rf_filter_coeff351_b(rf_filter_coeff351_b), 
		.rf_filter_coeff352_a(rf_filter_coeff352_a), 
		.rf_filter_coeff352_b(rf_filter_coeff352_b), 
		.rf_filter_coeff353_a(rf_filter_coeff353_a), 
		.rf_filter_coeff353_b(rf_filter_coeff353_b), 
		.rf_filter_coeff354_a(rf_filter_coeff354_a), 
		.rf_filter_coeff354_b(rf_filter_coeff354_b), 
		.rf_filter_coeff355_a(rf_filter_coeff355_a), 
		.rf_filter_coeff355_b(rf_filter_coeff355_b), 
		.rf_filter_coeff356_a(rf_filter_coeff356_a), 
		.rf_filter_coeff356_b(rf_filter_coeff356_b), 
		.rf_filter_coeff357_a(rf_filter_coeff357_a), 
		.rf_filter_coeff357_b(rf_filter_coeff357_b), 
		.rf_filter_coeff358_a(rf_filter_coeff358_a), 
		.rf_filter_coeff358_b(rf_filter_coeff358_b), 
		.rf_filter_coeff359_a(rf_filter_coeff359_a), 
		.rf_filter_coeff359_b(rf_filter_coeff359_b), 
		.rf_filter_coeff360_a(rf_filter_coeff360_a), 
		.rf_filter_coeff360_b(rf_filter_coeff360_b), 
		.rf_filter_coeff361_a(rf_filter_coeff361_a), 
		.rf_filter_coeff361_b(rf_filter_coeff361_b), 
		.rf_filter_coeff362_a(rf_filter_coeff362_a), 
		.rf_filter_coeff362_b(rf_filter_coeff362_b), 
		.rf_filter_coeff363_a(rf_filter_coeff363_a), 
		.rf_filter_coeff363_b(rf_filter_coeff363_b), 
		.rf_filter_coeff364_a(rf_filter_coeff364_a), 
		.rf_filter_coeff364_b(rf_filter_coeff364_b), 
		.rf_filter_coeff365_a(rf_filter_coeff365_a), 
		.rf_filter_coeff365_b(rf_filter_coeff365_b), 
		.rf_filter_coeff366_a(rf_filter_coeff366_a), 
		.rf_filter_coeff366_b(rf_filter_coeff366_b), 
		.rf_filter_coeff367_a(rf_filter_coeff367_a), 
		.rf_filter_coeff367_b(rf_filter_coeff367_b), 
		.rf_filter_coeff368_a(rf_filter_coeff368_a), 
		.rf_filter_coeff368_b(rf_filter_coeff368_b), 
		.rf_filter_coeff369_a(rf_filter_coeff369_a), 
		.rf_filter_coeff369_b(rf_filter_coeff369_b), 
		.rf_filter_coeff370_a(rf_filter_coeff370_a), 
		.rf_filter_coeff370_b(rf_filter_coeff370_b), 
		.rf_filter_coeff371_a(rf_filter_coeff371_a), 
		.rf_filter_coeff371_b(rf_filter_coeff371_b), 
		.rf_filter_coeff372_a(rf_filter_coeff372_a), 
		.rf_filter_coeff372_b(rf_filter_coeff372_b), 
		.rf_filter_coeff373_a(rf_filter_coeff373_a), 
		.rf_filter_coeff373_b(rf_filter_coeff373_b), 
		.rf_filter_coeff374_a(rf_filter_coeff374_a), 
		.rf_filter_coeff374_b(rf_filter_coeff374_b), 
		.rf_filter_coeff375_a(rf_filter_coeff375_a), 
		.rf_filter_coeff375_b(rf_filter_coeff375_b), 
		.rf_filter_coeff376_a(rf_filter_coeff376_a), 
		.rf_filter_coeff376_b(rf_filter_coeff376_b), 
		.rf_filter_coeff377_a(rf_filter_coeff377_a), 
		.rf_filter_coeff377_b(rf_filter_coeff377_b), 
		.rf_filter_coeff378_a(rf_filter_coeff378_a), 
		.rf_filter_coeff378_b(rf_filter_coeff378_b), 
		.rf_filter_coeff379_a(rf_filter_coeff379_a), 
		.rf_filter_coeff379_b(rf_filter_coeff379_b), 
		.rf_filter_coeff380_a(rf_filter_coeff380_a), 
		.rf_filter_coeff380_b(rf_filter_coeff380_b), 
		.rf_filter_coeff381_a(rf_filter_coeff381_a), 
		.rf_filter_coeff381_b(rf_filter_coeff381_b), 
		.rf_filter_coeff382_a(rf_filter_coeff382_a), 
		.rf_filter_coeff382_b(rf_filter_coeff382_b), 
		.rf_filter_coeff383_a(rf_filter_coeff383_a), 
		.rf_filter_coeff383_b(rf_filter_coeff383_b), 
		.rf_filter_coeff384_a(rf_filter_coeff384_a), 
		.rf_filter_coeff384_b(rf_filter_coeff384_b), 
		.rf_filter_coeff385_a(rf_filter_coeff385_a), 
		.rf_filter_coeff385_b(rf_filter_coeff385_b), 
		.rf_filter_coeff386_a(rf_filter_coeff386_a), 
		.rf_filter_coeff386_b(rf_filter_coeff386_b), 
		.rf_filter_coeff387_a(rf_filter_coeff387_a), 
		.rf_filter_coeff387_b(rf_filter_coeff387_b), 
		.rf_filter_coeff388_a(rf_filter_coeff388_a), 
		.rf_filter_coeff388_b(rf_filter_coeff388_b), 
		.rf_filter_coeff389_a(rf_filter_coeff389_a), 
		.rf_filter_coeff389_b(rf_filter_coeff389_b), 
		.rf_filter_coeff390_a(rf_filter_coeff390_a), 
		.rf_filter_coeff390_b(rf_filter_coeff390_b), 
		.rf_filter_coeff391_a(rf_filter_coeff391_a), 
		.rf_filter_coeff391_b(rf_filter_coeff391_b), 
		.rf_filter_coeff392_a(rf_filter_coeff392_a), 
		.rf_filter_coeff392_b(rf_filter_coeff392_b), 
		.rf_filter_coeff393_a(rf_filter_coeff393_a), 
		.rf_filter_coeff393_b(rf_filter_coeff393_b), 
		.rf_filter_coeff394_a(rf_filter_coeff394_a), 
		.rf_filter_coeff394_b(rf_filter_coeff394_b), 
		.rf_filter_coeff395_a(rf_filter_coeff395_a), 
		.rf_filter_coeff395_b(rf_filter_coeff395_b), 
		.rf_filter_coeff396_a(rf_filter_coeff396_a), 
		.rf_filter_coeff396_b(rf_filter_coeff396_b), 
		.rf_filter_coeff397_a(rf_filter_coeff397_a), 
		.rf_filter_coeff397_b(rf_filter_coeff397_b), 
		.rf_filter_coeff398_a(rf_filter_coeff398_a), 
		.rf_filter_coeff398_b(rf_filter_coeff398_b), 
		.rf_filter_coeff399_a(rf_filter_coeff399_a), 
		.rf_filter_coeff399_b(rf_filter_coeff399_b), 
		.rf_filter_coeff400_a(rf_filter_coeff400_a), 
		.rf_filter_coeff400_b(rf_filter_coeff400_b), 
		.rf_filter_coeff401_a(rf_filter_coeff401_a), 
		.rf_filter_coeff401_b(rf_filter_coeff401_b), 
		.rf_filter_coeff402_a(rf_filter_coeff402_a), 
		.rf_filter_coeff402_b(rf_filter_coeff402_b), 
		.rf_filter_coeff403_a(rf_filter_coeff403_a), 
		.rf_filter_coeff403_b(rf_filter_coeff403_b), 
		.rf_filter_coeff404_a(rf_filter_coeff404_a), 
		.rf_filter_coeff404_b(rf_filter_coeff404_b), 
		.rf_filter_coeff405_a(rf_filter_coeff405_a), 
		.rf_filter_coeff405_b(rf_filter_coeff405_b), 
		.rf_filter_coeff406_a(rf_filter_coeff406_a), 
		.rf_filter_coeff406_b(rf_filter_coeff406_b), 
		.rf_filter_coeff407_a(rf_filter_coeff407_a), 
		.rf_filter_coeff407_b(rf_filter_coeff407_b), 
		.rf_filter_coeff408_a(rf_filter_coeff408_a), 
		.rf_filter_coeff408_b(rf_filter_coeff408_b), 
		.rf_filter_coeff409_a(rf_filter_coeff409_a), 
		.rf_filter_coeff409_b(rf_filter_coeff409_b), 
		.rf_filter_coeff410_a(rf_filter_coeff410_a), 
		.rf_filter_coeff410_b(rf_filter_coeff410_b), 
		.rf_filter_coeff411_a(rf_filter_coeff411_a), 
		.rf_filter_coeff411_b(rf_filter_coeff411_b), 
		.rf_filter_coeff412_a(rf_filter_coeff412_a), 
		.rf_filter_coeff412_b(rf_filter_coeff412_b), 
		.rf_filter_coeff413_a(rf_filter_coeff413_a), 
		.rf_filter_coeff413_b(rf_filter_coeff413_b), 
		.rf_filter_coeff414_a(rf_filter_coeff414_a), 
		.rf_filter_coeff414_b(rf_filter_coeff414_b), 
		.rf_filter_coeff415_a(rf_filter_coeff415_a), 
		.rf_filter_coeff415_b(rf_filter_coeff415_b), 
		.rf_filter_coeff416_a(rf_filter_coeff416_a), 
		.rf_filter_coeff416_b(rf_filter_coeff416_b), 
		.rf_filter_coeff417_a(rf_filter_coeff417_a), 
		.rf_filter_coeff417_b(rf_filter_coeff417_b), 
		.rf_filter_coeff418_a(rf_filter_coeff418_a), 
		.rf_filter_coeff418_b(rf_filter_coeff418_b), 
		.rf_filter_coeff419_a(rf_filter_coeff419_a), 
		.rf_filter_coeff419_b(rf_filter_coeff419_b), 
		.rf_filter_coeff420_a(rf_filter_coeff420_a), 
		.rf_filter_coeff420_b(rf_filter_coeff420_b), 
		.rf_filter_coeff421_a(rf_filter_coeff421_a), 
		.rf_filter_coeff421_b(rf_filter_coeff421_b), 
		.rf_filter_coeff422_a(rf_filter_coeff422_a), 
		.rf_filter_coeff422_b(rf_filter_coeff422_b), 
		.rf_filter_coeff423_a(rf_filter_coeff423_a), 
		.rf_filter_coeff423_b(rf_filter_coeff423_b), 
		.rf_filter_coeff424_a(rf_filter_coeff424_a), 
		.rf_filter_coeff424_b(rf_filter_coeff424_b), 
		.rf_filter_coeff425_a(rf_filter_coeff425_a), 
		.rf_filter_coeff425_b(rf_filter_coeff425_b), 
		.rf_filter_coeff426_a(rf_filter_coeff426_a), 
		.rf_filter_coeff426_b(rf_filter_coeff426_b), 
		.rf_filter_coeff427_a(rf_filter_coeff427_a), 
		.rf_filter_coeff427_b(rf_filter_coeff427_b), 
		.rf_filter_coeff428_a(rf_filter_coeff428_a), 
		.rf_filter_coeff428_b(rf_filter_coeff428_b), 
		.rf_filter_coeff429_a(rf_filter_coeff429_a), 
		.rf_filter_coeff429_b(rf_filter_coeff429_b), 
		.rf_filter_coeff430_a(rf_filter_coeff430_a), 
		.rf_filter_coeff430_b(rf_filter_coeff430_b), 
		.rf_filter_coeff431_a(rf_filter_coeff431_a), 
		.rf_filter_coeff431_b(rf_filter_coeff431_b), 
		.rf_filter_coeff432_a(rf_filter_coeff432_a), 
		.rf_filter_coeff432_b(rf_filter_coeff432_b), 
		.rf_filter_coeff433_a(rf_filter_coeff433_a), 
		.rf_filter_coeff433_b(rf_filter_coeff433_b), 
		.rf_filter_coeff434_a(rf_filter_coeff434_a), 
		.rf_filter_coeff434_b(rf_filter_coeff434_b), 
		.rf_filter_coeff435_a(rf_filter_coeff435_a), 
		.rf_filter_coeff435_b(rf_filter_coeff435_b), 
		.rf_filter_coeff436_a(rf_filter_coeff436_a), 
		.rf_filter_coeff436_b(rf_filter_coeff436_b), 
		.rf_filter_coeff437_a(rf_filter_coeff437_a), 
		.rf_filter_coeff437_b(rf_filter_coeff437_b), 
		.rf_filter_coeff438_a(rf_filter_coeff438_a), 
		.rf_filter_coeff438_b(rf_filter_coeff438_b), 
		.rf_filter_coeff439_a(rf_filter_coeff439_a), 
		.rf_filter_coeff439_b(rf_filter_coeff439_b), 
		.rf_filter_coeff440_a(rf_filter_coeff440_a), 
		.rf_filter_coeff440_b(rf_filter_coeff440_b), 
		.rf_filter_coeff441_a(rf_filter_coeff441_a), 
		.rf_filter_coeff441_b(rf_filter_coeff441_b), 
		.rf_filter_coeff442_a(rf_filter_coeff442_a), 
		.rf_filter_coeff442_b(rf_filter_coeff442_b), 
		.rf_filter_coeff443_a(rf_filter_coeff443_a), 
		.rf_filter_coeff443_b(rf_filter_coeff443_b), 
		.rf_filter_coeff444_a(rf_filter_coeff444_a), 
		.rf_filter_coeff444_b(rf_filter_coeff444_b), 
		.rf_filter_coeff445_a(rf_filter_coeff445_a), 
		.rf_filter_coeff445_b(rf_filter_coeff445_b), 
		.rf_filter_coeff446_a(rf_filter_coeff446_a), 
		.rf_filter_coeff446_b(rf_filter_coeff446_b), 
		.rf_filter_coeff447_a(rf_filter_coeff447_a), 
		.rf_filter_coeff447_b(rf_filter_coeff447_b), 
		.rf_filter_coeff448_a(rf_filter_coeff448_a), 
		.rf_filter_coeff448_b(rf_filter_coeff448_b), 
		.rf_filter_coeff449_a(rf_filter_coeff449_a), 
		.rf_filter_coeff449_b(rf_filter_coeff449_b), 
		.rf_filter_coeff450_a(rf_filter_coeff450_a), 
		.rf_filter_coeff450_b(rf_filter_coeff450_b), 
		.rf_filter_coeff451_a(rf_filter_coeff451_a), 
		.rf_filter_coeff451_b(rf_filter_coeff451_b), 
		.rf_filter_coeff452_a(rf_filter_coeff452_a), 
		.rf_filter_coeff452_b(rf_filter_coeff452_b), 
		.rf_filter_coeff453_a(rf_filter_coeff453_a), 
		.rf_filter_coeff453_b(rf_filter_coeff453_b), 
		.rf_filter_coeff454_a(rf_filter_coeff454_a), 
		.rf_filter_coeff454_b(rf_filter_coeff454_b), 
		.rf_filter_coeff455_a(rf_filter_coeff455_a), 
		.rf_filter_coeff455_b(rf_filter_coeff455_b), 
		.rf_filter_coeff456_a(rf_filter_coeff456_a), 
		.rf_filter_coeff456_b(rf_filter_coeff456_b), 
		.rf_filter_coeff457_a(rf_filter_coeff457_a), 
		.rf_filter_coeff457_b(rf_filter_coeff457_b), 
		.rf_filter_coeff458_a(rf_filter_coeff458_a), 
		.rf_filter_coeff458_b(rf_filter_coeff458_b), 
		.rf_filter_coeff459_a(rf_filter_coeff459_a), 
		.rf_filter_coeff459_b(rf_filter_coeff459_b), 
		.rf_filter_coeff460_a(rf_filter_coeff460_a), 
		.rf_filter_coeff460_b(rf_filter_coeff460_b), 
		.rf_filter_coeff461_a(rf_filter_coeff461_a), 
		.rf_filter_coeff461_b(rf_filter_coeff461_b), 
		.rf_filter_coeff462_a(rf_filter_coeff462_a), 
		.rf_filter_coeff462_b(rf_filter_coeff462_b), 
		.rf_filter_coeff463_a(rf_filter_coeff463_a), 
		.rf_filter_coeff463_b(rf_filter_coeff463_b), 
		.rf_filter_coeff464_a(rf_filter_coeff464_a), 
		.rf_filter_coeff464_b(rf_filter_coeff464_b), 
		.rf_filter_coeff465_a(rf_filter_coeff465_a), 
		.rf_filter_coeff465_b(rf_filter_coeff465_b), 
		.rf_filter_coeff466_a(rf_filter_coeff466_a), 
		.rf_filter_coeff466_b(rf_filter_coeff466_b), 
		.rf_filter_coeff467_a(rf_filter_coeff467_a), 
		.rf_filter_coeff467_b(rf_filter_coeff467_b), 
		.rf_filter_coeff468_a(rf_filter_coeff468_a), 
		.rf_filter_coeff468_b(rf_filter_coeff468_b), 
		.rf_filter_coeff469_a(rf_filter_coeff469_a), 
		.rf_filter_coeff469_b(rf_filter_coeff469_b), 
		.rf_filter_coeff470_a(rf_filter_coeff470_a), 
		.rf_filter_coeff470_b(rf_filter_coeff470_b), 
		.rf_filter_coeff471_a(rf_filter_coeff471_a), 
		.rf_filter_coeff471_b(rf_filter_coeff471_b), 
		.rf_filter_coeff472_a(rf_filter_coeff472_a), 
		.rf_filter_coeff472_b(rf_filter_coeff472_b), 
		.rf_filter_coeff473_a(rf_filter_coeff473_a), 
		.rf_filter_coeff473_b(rf_filter_coeff473_b), 
		.rf_filter_coeff474_a(rf_filter_coeff474_a), 
		.rf_filter_coeff474_b(rf_filter_coeff474_b), 
		.rf_filter_coeff475_a(rf_filter_coeff475_a), 
		.rf_filter_coeff475_b(rf_filter_coeff475_b), 
		.rf_filter_coeff476_a(rf_filter_coeff476_a), 
		.rf_filter_coeff476_b(rf_filter_coeff476_b), 
		.rf_filter_coeff477_a(rf_filter_coeff477_a), 
		.rf_filter_coeff477_b(rf_filter_coeff477_b), 
		.rf_filter_coeff478_a(rf_filter_coeff478_a), 
		.rf_filter_coeff478_b(rf_filter_coeff478_b), 
		.rf_filter_coeff479_a(rf_filter_coeff479_a), 
		.rf_filter_coeff479_b(rf_filter_coeff479_b), 
		.rf_filter_coeff480_a(rf_filter_coeff480_a), 
		.rf_filter_coeff480_b(rf_filter_coeff480_b), 
		.rf_filter_coeff481_a(rf_filter_coeff481_a), 
		.rf_filter_coeff481_b(rf_filter_coeff481_b), 
		.rf_filter_coeff482_a(rf_filter_coeff482_a), 
		.rf_filter_coeff482_b(rf_filter_coeff482_b), 
		.rf_filter_coeff483_a(rf_filter_coeff483_a), 
		.rf_filter_coeff483_b(rf_filter_coeff483_b), 
		.rf_filter_coeff484_a(rf_filter_coeff484_a), 
		.rf_filter_coeff484_b(rf_filter_coeff484_b), 
		.rf_filter_coeff485_a(rf_filter_coeff485_a), 
		.rf_filter_coeff485_b(rf_filter_coeff485_b), 
		.rf_filter_coeff486_a(rf_filter_coeff486_a), 
		.rf_filter_coeff486_b(rf_filter_coeff486_b), 
		.rf_filter_coeff487_a(rf_filter_coeff487_a), 
		.rf_filter_coeff487_b(rf_filter_coeff487_b), 
		.rf_filter_coeff488_a(rf_filter_coeff488_a), 
		.rf_filter_coeff488_b(rf_filter_coeff488_b), 
		.rf_filter_coeff489_a(rf_filter_coeff489_a), 
		.rf_filter_coeff489_b(rf_filter_coeff489_b), 
		.rf_filter_coeff490_a(rf_filter_coeff490_a), 
		.rf_filter_coeff490_b(rf_filter_coeff490_b), 
		.rf_filter_coeff491_a(rf_filter_coeff491_a), 
		.rf_filter_coeff491_b(rf_filter_coeff491_b), 
		.rf_filter_coeff492_a(rf_filter_coeff492_a), 
		.rf_filter_coeff492_b(rf_filter_coeff492_b), 
		.rf_filter_coeff493_a(rf_filter_coeff493_a), 
		.rf_filter_coeff493_b(rf_filter_coeff493_b), 
		.rf_filter_coeff494_a(rf_filter_coeff494_a), 
		.rf_filter_coeff494_b(rf_filter_coeff494_b), 
		.rf_filter_coeff495_a(rf_filter_coeff495_a), 
		.rf_filter_coeff495_b(rf_filter_coeff495_b), 
		.rf_filter_coeff496_a(rf_filter_coeff496_a), 
		.rf_filter_coeff496_b(rf_filter_coeff496_b), 
		.rf_filter_coeff497_a(rf_filter_coeff497_a), 
		.rf_filter_coeff497_b(rf_filter_coeff497_b), 
		.rf_filter_coeff498_a(rf_filter_coeff498_a), 
		.rf_filter_coeff498_b(rf_filter_coeff498_b), 
		.rf_filter_coeff499_a(rf_filter_coeff499_a), 
		.rf_filter_coeff499_b(rf_filter_coeff499_b), 
		.rf_filter_coeff500_a(rf_filter_coeff500_a), 
		.rf_filter_coeff500_b(rf_filter_coeff500_b), 
		.rf_filter_coeff501_a(rf_filter_coeff501_a), 
		.rf_filter_coeff501_b(rf_filter_coeff501_b), 
		.rf_filter_coeff502_a(rf_filter_coeff502_a), 
		.rf_filter_coeff502_b(rf_filter_coeff502_b), 
		.rf_filter_coeff503_a(rf_filter_coeff503_a), 
		.rf_filter_coeff503_b(rf_filter_coeff503_b), 
		.rf_filter_coeff504_a(rf_filter_coeff504_a), 
		.rf_filter_coeff504_b(rf_filter_coeff504_b), 
		.rf_filter_coeff505_a(rf_filter_coeff505_a), 
		.rf_filter_coeff505_b(rf_filter_coeff505_b), 
		.rf_filter_coeff506_a(rf_filter_coeff506_a), 
		.rf_filter_coeff506_b(rf_filter_coeff506_b), 
		.rf_filter_coeff507_a(rf_filter_coeff507_a), 
		.rf_filter_coeff507_b(rf_filter_coeff507_b), 
		.rf_filter_coeff508_a(rf_filter_coeff508_a), 
		.rf_filter_coeff508_b(rf_filter_coeff508_b), 
		.rf_filter_coeff509_a(rf_filter_coeff509_a), 
		.rf_filter_coeff509_b(rf_filter_coeff509_b), 
		.rf_filter_coeff510_a(rf_filter_coeff510_a), 
		.rf_filter_coeff510_b(rf_filter_coeff510_b), 
		.rf_filter_coeff511_a(rf_filter_coeff511_a), 
		.rf_filter_coeff511_b(rf_filter_coeff511_b)
	);

	initial begin
		// Initialize Inputs
		rst_n = 0;
		clk = 0;
		addr = 0;
		wdata = 0;
		w_enable = 0;
		wxfc = 0;
		ro_fifo_underrun = 0;
		ro_fifo_overrun = 0;
		ro_filter_ovf_flag = 0;

		// Wait 100 ns for global reset to finish
		#100;
		
		
	end
	
      
endmodule

