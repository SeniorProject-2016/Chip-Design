`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:31:00 02/09/2016
// Design Name:   filter
// Module Name:   Z:/Desktop/chip/filter_tf_test_xfc.v
// Project Name:  chip
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: filter
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module filter_tf_test_xfc;

	// Inputs
	reg clk;
	reg rstb;
	reg [31:0] filt_input_data;
	reg aud_in_rts;
	reg aud_out_rtr;
	reg [2:0] rf_filter_shift;
	reg rf_filter_clip_en;
	reg trig_filter_ovf_flag_clear;
	reg [7:0] rf_filter_coeff0_a;
	reg [7:0] rf_filter_coeff0_b;
	reg [7:0] rf_filter_coeff1_a;
	reg [7:0] rf_filter_coeff1_b;
	reg [7:0] rf_filter_coeff2_a;
	reg [7:0] rf_filter_coeff2_b;
	reg [7:0] rf_filter_coeff3_a;
	reg [7:0] rf_filter_coeff3_b;
	reg [7:0] rf_filter_coeff4_a;
	reg [7:0] rf_filter_coeff4_b;
	reg [7:0] rf_filter_coeff5_a;
	reg [7:0] rf_filter_coeff5_b;
	reg [7:0] rf_filter_coeff6_a;
	reg [7:0] rf_filter_coeff6_b;
	reg [7:0] rf_filter_coeff7_a;
	reg [7:0] rf_filter_coeff7_b;
	reg [7:0] rf_filter_coeff8_a;
	reg [7:0] rf_filter_coeff8_b;
	reg [7:0] rf_filter_coeff9_a;
	reg [7:0] rf_filter_coeff9_b;
	reg [7:0] rf_filter_coeff10_a;
	reg [7:0] rf_filter_coeff10_b;
	reg [7:0] rf_filter_coeff11_a;
	reg [7:0] rf_filter_coeff11_b;
	reg [7:0] rf_filter_coeff12_a;
	reg [7:0] rf_filter_coeff12_b;
	reg [7:0] rf_filter_coeff13_a;
	reg [7:0] rf_filter_coeff13_b;
	reg [7:0] rf_filter_coeff14_a;
	reg [7:0] rf_filter_coeff14_b;
	reg [7:0] rf_filter_coeff15_a;
	reg [7:0] rf_filter_coeff15_b;
	reg [7:0] rf_filter_coeff16_a;
	reg [7:0] rf_filter_coeff16_b;
	reg [7:0] rf_filter_coeff17_a;
	reg [7:0] rf_filter_coeff17_b;
	reg [7:0] rf_filter_coeff18_a;
	reg [7:0] rf_filter_coeff18_b;
	reg [7:0] rf_filter_coeff19_a;
	reg [7:0] rf_filter_coeff19_b;
	reg [7:0] rf_filter_coeff20_a;
	reg [7:0] rf_filter_coeff20_b;
	reg [7:0] rf_filter_coeff21_a;
	reg [7:0] rf_filter_coeff21_b;
	reg [7:0] rf_filter_coeff22_a;
	reg [7:0] rf_filter_coeff22_b;
	reg [7:0] rf_filter_coeff23_a;
	reg [7:0] rf_filter_coeff23_b;
	reg [7:0] rf_filter_coeff24_a;
	reg [7:0] rf_filter_coeff24_b;
	reg [7:0] rf_filter_coeff25_a;
	reg [7:0] rf_filter_coeff25_b;
	reg [7:0] rf_filter_coeff26_a;
	reg [7:0] rf_filter_coeff26_b;
	reg [7:0] rf_filter_coeff27_a;
	reg [7:0] rf_filter_coeff27_b;
	reg [7:0] rf_filter_coeff28_a;
	reg [7:0] rf_filter_coeff28_b;
	reg [7:0] rf_filter_coeff29_a;
	reg [7:0] rf_filter_coeff29_b;
	reg [7:0] rf_filter_coeff30_a;
	reg [7:0] rf_filter_coeff30_b;
	reg [7:0] rf_filter_coeff31_a;
	reg [7:0] rf_filter_coeff31_b;
	reg [7:0] rf_filter_coeff32_a;
	reg [7:0] rf_filter_coeff32_b;
	reg [7:0] rf_filter_coeff33_a;
	reg [7:0] rf_filter_coeff33_b;
	reg [7:0] rf_filter_coeff34_a;
	reg [7:0] rf_filter_coeff34_b;
	reg [7:0] rf_filter_coeff35_a;
	reg [7:0] rf_filter_coeff35_b;
	reg [7:0] rf_filter_coeff36_a;
	reg [7:0] rf_filter_coeff36_b;
	reg [7:0] rf_filter_coeff37_a;
	reg [7:0] rf_filter_coeff37_b;
	reg [7:0] rf_filter_coeff38_a;
	reg [7:0] rf_filter_coeff38_b;
	reg [7:0] rf_filter_coeff39_a;
	reg [7:0] rf_filter_coeff39_b;
	reg [7:0] rf_filter_coeff40_a;
	reg [7:0] rf_filter_coeff40_b;
	reg [7:0] rf_filter_coeff41_a;
	reg [7:0] rf_filter_coeff41_b;
	reg [7:0] rf_filter_coeff42_a;
	reg [7:0] rf_filter_coeff42_b;
	reg [7:0] rf_filter_coeff43_a;
	reg [7:0] rf_filter_coeff43_b;
	reg [7:0] rf_filter_coeff44_a;
	reg [7:0] rf_filter_coeff44_b;
	reg [7:0] rf_filter_coeff45_a;
	reg [7:0] rf_filter_coeff45_b;
	reg [7:0] rf_filter_coeff46_a;
	reg [7:0] rf_filter_coeff46_b;
	reg [7:0] rf_filter_coeff47_a;
	reg [7:0] rf_filter_coeff47_b;
	reg [7:0] rf_filter_coeff48_a;
	reg [7:0] rf_filter_coeff48_b;
	reg [7:0] rf_filter_coeff49_a;
	reg [7:0] rf_filter_coeff49_b;
	reg [7:0] rf_filter_coeff50_a;
	reg [7:0] rf_filter_coeff50_b;
	reg [7:0] rf_filter_coeff51_a;
	reg [7:0] rf_filter_coeff51_b;
	reg [7:0] rf_filter_coeff52_a;
	reg [7:0] rf_filter_coeff52_b;
	reg [7:0] rf_filter_coeff53_a;
	reg [7:0] rf_filter_coeff53_b;
	reg [7:0] rf_filter_coeff54_a;
	reg [7:0] rf_filter_coeff54_b;
	reg [7:0] rf_filter_coeff55_a;
	reg [7:0] rf_filter_coeff55_b;
	reg [7:0] rf_filter_coeff56_a;
	reg [7:0] rf_filter_coeff56_b;
	reg [7:0] rf_filter_coeff57_a;
	reg [7:0] rf_filter_coeff57_b;
	reg [7:0] rf_filter_coeff58_a;
	reg [7:0] rf_filter_coeff58_b;
	reg [7:0] rf_filter_coeff59_a;
	reg [7:0] rf_filter_coeff59_b;
	reg [7:0] rf_filter_coeff60_a;
	reg [7:0] rf_filter_coeff60_b;
	reg [7:0] rf_filter_coeff61_a;
	reg [7:0] rf_filter_coeff61_b;
	reg [7:0] rf_filter_coeff62_a;
	reg [7:0] rf_filter_coeff62_b;
	reg [7:0] rf_filter_coeff63_a;
	reg [7:0] rf_filter_coeff63_b;
	reg [7:0] rf_filter_coeff64_a;
	reg [7:0] rf_filter_coeff64_b;
	reg [7:0] rf_filter_coeff65_a;
	reg [7:0] rf_filter_coeff65_b;
	reg [7:0] rf_filter_coeff66_a;
	reg [7:0] rf_filter_coeff66_b;
	reg [7:0] rf_filter_coeff67_a;
	reg [7:0] rf_filter_coeff67_b;
	reg [7:0] rf_filter_coeff68_a;
	reg [7:0] rf_filter_coeff68_b;
	reg [7:0] rf_filter_coeff69_a;
	reg [7:0] rf_filter_coeff69_b;
	reg [7:0] rf_filter_coeff70_a;
	reg [7:0] rf_filter_coeff70_b;
	reg [7:0] rf_filter_coeff71_a;
	reg [7:0] rf_filter_coeff71_b;
	reg [7:0] rf_filter_coeff72_a;
	reg [7:0] rf_filter_coeff72_b;
	reg [7:0] rf_filter_coeff73_a;
	reg [7:0] rf_filter_coeff73_b;
	reg [7:0] rf_filter_coeff74_a;
	reg [7:0] rf_filter_coeff74_b;
	reg [7:0] rf_filter_coeff75_a;
	reg [7:0] rf_filter_coeff75_b;
	reg [7:0] rf_filter_coeff76_a;
	reg [7:0] rf_filter_coeff76_b;
	reg [7:0] rf_filter_coeff77_a;
	reg [7:0] rf_filter_coeff77_b;
	reg [7:0] rf_filter_coeff78_a;
	reg [7:0] rf_filter_coeff78_b;
	reg [7:0] rf_filter_coeff79_a;
	reg [7:0] rf_filter_coeff79_b;
	reg [7:0] rf_filter_coeff80_a;
	reg [7:0] rf_filter_coeff80_b;
	reg [7:0] rf_filter_coeff81_a;
	reg [7:0] rf_filter_coeff81_b;
	reg [7:0] rf_filter_coeff82_a;
	reg [7:0] rf_filter_coeff82_b;
	reg [7:0] rf_filter_coeff83_a;
	reg [7:0] rf_filter_coeff83_b;
	reg [7:0] rf_filter_coeff84_a;
	reg [7:0] rf_filter_coeff84_b;
	reg [7:0] rf_filter_coeff85_a;
	reg [7:0] rf_filter_coeff85_b;
	reg [7:0] rf_filter_coeff86_a;
	reg [7:0] rf_filter_coeff86_b;
	reg [7:0] rf_filter_coeff87_a;
	reg [7:0] rf_filter_coeff87_b;
	reg [7:0] rf_filter_coeff88_a;
	reg [7:0] rf_filter_coeff88_b;
	reg [7:0] rf_filter_coeff89_a;
	reg [7:0] rf_filter_coeff89_b;
	reg [7:0] rf_filter_coeff90_a;
	reg [7:0] rf_filter_coeff90_b;
	reg [7:0] rf_filter_coeff91_a;
	reg [7:0] rf_filter_coeff91_b;
	reg [7:0] rf_filter_coeff92_a;
	reg [7:0] rf_filter_coeff92_b;
	reg [7:0] rf_filter_coeff93_a;
	reg [7:0] rf_filter_coeff93_b;
	reg [7:0] rf_filter_coeff94_a;
	reg [7:0] rf_filter_coeff94_b;
	reg [7:0] rf_filter_coeff95_a;
	reg [7:0] rf_filter_coeff95_b;
	reg [7:0] rf_filter_coeff96_a;
	reg [7:0] rf_filter_coeff96_b;
	reg [7:0] rf_filter_coeff97_a;
	reg [7:0] rf_filter_coeff97_b;
	reg [7:0] rf_filter_coeff98_a;
	reg [7:0] rf_filter_coeff98_b;
	reg [7:0] rf_filter_coeff99_a;
	reg [7:0] rf_filter_coeff99_b;
	reg [7:0] rf_filter_coeff100_a;
	reg [7:0] rf_filter_coeff100_b;
	reg [7:0] rf_filter_coeff101_a;
	reg [7:0] rf_filter_coeff101_b;
	reg [7:0] rf_filter_coeff102_a;
	reg [7:0] rf_filter_coeff102_b;
	reg [7:0] rf_filter_coeff103_a;
	reg [7:0] rf_filter_coeff103_b;
	reg [7:0] rf_filter_coeff104_a;
	reg [7:0] rf_filter_coeff104_b;
	reg [7:0] rf_filter_coeff105_a;
	reg [7:0] rf_filter_coeff105_b;
	reg [7:0] rf_filter_coeff106_a;
	reg [7:0] rf_filter_coeff106_b;
	reg [7:0] rf_filter_coeff107_a;
	reg [7:0] rf_filter_coeff107_b;
	reg [7:0] rf_filter_coeff108_a;
	reg [7:0] rf_filter_coeff108_b;
	reg [7:0] rf_filter_coeff109_a;
	reg [7:0] rf_filter_coeff109_b;
	reg [7:0] rf_filter_coeff110_a;
	reg [7:0] rf_filter_coeff110_b;
	reg [7:0] rf_filter_coeff111_a;
	reg [7:0] rf_filter_coeff111_b;
	reg [7:0] rf_filter_coeff112_a;
	reg [7:0] rf_filter_coeff112_b;
	reg [7:0] rf_filter_coeff113_a;
	reg [7:0] rf_filter_coeff113_b;
	reg [7:0] rf_filter_coeff114_a;
	reg [7:0] rf_filter_coeff114_b;
	reg [7:0] rf_filter_coeff115_a;
	reg [7:0] rf_filter_coeff115_b;
	reg [7:0] rf_filter_coeff116_a;
	reg [7:0] rf_filter_coeff116_b;
	reg [7:0] rf_filter_coeff117_a;
	reg [7:0] rf_filter_coeff117_b;
	reg [7:0] rf_filter_coeff118_a;
	reg [7:0] rf_filter_coeff118_b;
	reg [7:0] rf_filter_coeff119_a;
	reg [7:0] rf_filter_coeff119_b;
	reg [7:0] rf_filter_coeff120_a;
	reg [7:0] rf_filter_coeff120_b;
	reg [7:0] rf_filter_coeff121_a;
	reg [7:0] rf_filter_coeff121_b;
	reg [7:0] rf_filter_coeff122_a;
	reg [7:0] rf_filter_coeff122_b;
	reg [7:0] rf_filter_coeff123_a;
	reg [7:0] rf_filter_coeff123_b;
	reg [7:0] rf_filter_coeff124_a;
	reg [7:0] rf_filter_coeff124_b;
	reg [7:0] rf_filter_coeff125_a;
	reg [7:0] rf_filter_coeff125_b;
	reg [7:0] rf_filter_coeff126_a;
	reg [7:0] rf_filter_coeff126_b;
	reg [7:0] rf_filter_coeff127_a;
	reg [7:0] rf_filter_coeff127_b;
	reg [7:0] rf_filter_coeff128_a;
	reg [7:0] rf_filter_coeff128_b;
	reg [7:0] rf_filter_coeff129_a;
	reg [7:0] rf_filter_coeff129_b;
	reg [7:0] rf_filter_coeff130_a;
	reg [7:0] rf_filter_coeff130_b;
	reg [7:0] rf_filter_coeff131_a;
	reg [7:0] rf_filter_coeff131_b;
	reg [7:0] rf_filter_coeff132_a;
	reg [7:0] rf_filter_coeff132_b;
	reg [7:0] rf_filter_coeff133_a;
	reg [7:0] rf_filter_coeff133_b;
	reg [7:0] rf_filter_coeff134_a;
	reg [7:0] rf_filter_coeff134_b;
	reg [7:0] rf_filter_coeff135_a;
	reg [7:0] rf_filter_coeff135_b;
	reg [7:0] rf_filter_coeff136_a;
	reg [7:0] rf_filter_coeff136_b;
	reg [7:0] rf_filter_coeff137_a;
	reg [7:0] rf_filter_coeff137_b;
	reg [7:0] rf_filter_coeff138_a;
	reg [7:0] rf_filter_coeff138_b;
	reg [7:0] rf_filter_coeff139_a;
	reg [7:0] rf_filter_coeff139_b;
	reg [7:0] rf_filter_coeff140_a;
	reg [7:0] rf_filter_coeff140_b;
	reg [7:0] rf_filter_coeff141_a;
	reg [7:0] rf_filter_coeff141_b;
	reg [7:0] rf_filter_coeff142_a;
	reg [7:0] rf_filter_coeff142_b;
	reg [7:0] rf_filter_coeff143_a;
	reg [7:0] rf_filter_coeff143_b;
	reg [7:0] rf_filter_coeff144_a;
	reg [7:0] rf_filter_coeff144_b;
	reg [7:0] rf_filter_coeff145_a;
	reg [7:0] rf_filter_coeff145_b;
	reg [7:0] rf_filter_coeff146_a;
	reg [7:0] rf_filter_coeff146_b;
	reg [7:0] rf_filter_coeff147_a;
	reg [7:0] rf_filter_coeff147_b;
	reg [7:0] rf_filter_coeff148_a;
	reg [7:0] rf_filter_coeff148_b;
	reg [7:0] rf_filter_coeff149_a;
	reg [7:0] rf_filter_coeff149_b;
	reg [7:0] rf_filter_coeff150_a;
	reg [7:0] rf_filter_coeff150_b;
	reg [7:0] rf_filter_coeff151_a;
	reg [7:0] rf_filter_coeff151_b;
	reg [7:0] rf_filter_coeff152_a;
	reg [7:0] rf_filter_coeff152_b;
	reg [7:0] rf_filter_coeff153_a;
	reg [7:0] rf_filter_coeff153_b;
	reg [7:0] rf_filter_coeff154_a;
	reg [7:0] rf_filter_coeff154_b;
	reg [7:0] rf_filter_coeff155_a;
	reg [7:0] rf_filter_coeff155_b;
	reg [7:0] rf_filter_coeff156_a;
	reg [7:0] rf_filter_coeff156_b;
	reg [7:0] rf_filter_coeff157_a;
	reg [7:0] rf_filter_coeff157_b;
	reg [7:0] rf_filter_coeff158_a;
	reg [7:0] rf_filter_coeff158_b;
	reg [7:0] rf_filter_coeff159_a;
	reg [7:0] rf_filter_coeff159_b;
	reg [7:0] rf_filter_coeff160_a;
	reg [7:0] rf_filter_coeff160_b;
	reg [7:0] rf_filter_coeff161_a;
	reg [7:0] rf_filter_coeff161_b;
	reg [7:0] rf_filter_coeff162_a;
	reg [7:0] rf_filter_coeff162_b;
	reg [7:0] rf_filter_coeff163_a;
	reg [7:0] rf_filter_coeff163_b;
	reg [7:0] rf_filter_coeff164_a;
	reg [7:0] rf_filter_coeff164_b;
	reg [7:0] rf_filter_coeff165_a;
	reg [7:0] rf_filter_coeff165_b;
	reg [7:0] rf_filter_coeff166_a;
	reg [7:0] rf_filter_coeff166_b;
	reg [7:0] rf_filter_coeff167_a;
	reg [7:0] rf_filter_coeff167_b;
	reg [7:0] rf_filter_coeff168_a;
	reg [7:0] rf_filter_coeff168_b;
	reg [7:0] rf_filter_coeff169_a;
	reg [7:0] rf_filter_coeff169_b;
	reg [7:0] rf_filter_coeff170_a;
	reg [7:0] rf_filter_coeff170_b;
	reg [7:0] rf_filter_coeff171_a;
	reg [7:0] rf_filter_coeff171_b;
	reg [7:0] rf_filter_coeff172_a;
	reg [7:0] rf_filter_coeff172_b;
	reg [7:0] rf_filter_coeff173_a;
	reg [7:0] rf_filter_coeff173_b;
	reg [7:0] rf_filter_coeff174_a;
	reg [7:0] rf_filter_coeff174_b;
	reg [7:0] rf_filter_coeff175_a;
	reg [7:0] rf_filter_coeff175_b;
	reg [7:0] rf_filter_coeff176_a;
	reg [7:0] rf_filter_coeff176_b;
	reg [7:0] rf_filter_coeff177_a;
	reg [7:0] rf_filter_coeff177_b;
	reg [7:0] rf_filter_coeff178_a;
	reg [7:0] rf_filter_coeff178_b;
	reg [7:0] rf_filter_coeff179_a;
	reg [7:0] rf_filter_coeff179_b;
	reg [7:0] rf_filter_coeff180_a;
	reg [7:0] rf_filter_coeff180_b;
	reg [7:0] rf_filter_coeff181_a;
	reg [7:0] rf_filter_coeff181_b;
	reg [7:0] rf_filter_coeff182_a;
	reg [7:0] rf_filter_coeff182_b;
	reg [7:0] rf_filter_coeff183_a;
	reg [7:0] rf_filter_coeff183_b;
	reg [7:0] rf_filter_coeff184_a;
	reg [7:0] rf_filter_coeff184_b;
	reg [7:0] rf_filter_coeff185_a;
	reg [7:0] rf_filter_coeff185_b;
	reg [7:0] rf_filter_coeff186_a;
	reg [7:0] rf_filter_coeff186_b;
	reg [7:0] rf_filter_coeff187_a;
	reg [7:0] rf_filter_coeff187_b;
	reg [7:0] rf_filter_coeff188_a;
	reg [7:0] rf_filter_coeff188_b;
	reg [7:0] rf_filter_coeff189_a;
	reg [7:0] rf_filter_coeff189_b;
	reg [7:0] rf_filter_coeff190_a;
	reg [7:0] rf_filter_coeff190_b;
	reg [7:0] rf_filter_coeff191_a;
	reg [7:0] rf_filter_coeff191_b;
	reg [7:0] rf_filter_coeff192_a;
	reg [7:0] rf_filter_coeff192_b;
	reg [7:0] rf_filter_coeff193_a;
	reg [7:0] rf_filter_coeff193_b;
	reg [7:0] rf_filter_coeff194_a;
	reg [7:0] rf_filter_coeff194_b;
	reg [7:0] rf_filter_coeff195_a;
	reg [7:0] rf_filter_coeff195_b;
	reg [7:0] rf_filter_coeff196_a;
	reg [7:0] rf_filter_coeff196_b;
	reg [7:0] rf_filter_coeff197_a;
	reg [7:0] rf_filter_coeff197_b;
	reg [7:0] rf_filter_coeff198_a;
	reg [7:0] rf_filter_coeff198_b;
	reg [7:0] rf_filter_coeff199_a;
	reg [7:0] rf_filter_coeff199_b;
	reg [7:0] rf_filter_coeff200_a;
	reg [7:0] rf_filter_coeff200_b;
	reg [7:0] rf_filter_coeff201_a;
	reg [7:0] rf_filter_coeff201_b;
	reg [7:0] rf_filter_coeff202_a;
	reg [7:0] rf_filter_coeff202_b;
	reg [7:0] rf_filter_coeff203_a;
	reg [7:0] rf_filter_coeff203_b;
	reg [7:0] rf_filter_coeff204_a;
	reg [7:0] rf_filter_coeff204_b;
	reg [7:0] rf_filter_coeff205_a;
	reg [7:0] rf_filter_coeff205_b;
	reg [7:0] rf_filter_coeff206_a;
	reg [7:0] rf_filter_coeff206_b;
	reg [7:0] rf_filter_coeff207_a;
	reg [7:0] rf_filter_coeff207_b;
	reg [7:0] rf_filter_coeff208_a;
	reg [7:0] rf_filter_coeff208_b;
	reg [7:0] rf_filter_coeff209_a;
	reg [7:0] rf_filter_coeff209_b;
	reg [7:0] rf_filter_coeff210_a;
	reg [7:0] rf_filter_coeff210_b;
	reg [7:0] rf_filter_coeff211_a;
	reg [7:0] rf_filter_coeff211_b;
	reg [7:0] rf_filter_coeff212_a;
	reg [7:0] rf_filter_coeff212_b;
	reg [7:0] rf_filter_coeff213_a;
	reg [7:0] rf_filter_coeff213_b;
	reg [7:0] rf_filter_coeff214_a;
	reg [7:0] rf_filter_coeff214_b;
	reg [7:0] rf_filter_coeff215_a;
	reg [7:0] rf_filter_coeff215_b;
	reg [7:0] rf_filter_coeff216_a;
	reg [7:0] rf_filter_coeff216_b;
	reg [7:0] rf_filter_coeff217_a;
	reg [7:0] rf_filter_coeff217_b;
	reg [7:0] rf_filter_coeff218_a;
	reg [7:0] rf_filter_coeff218_b;
	reg [7:0] rf_filter_coeff219_a;
	reg [7:0] rf_filter_coeff219_b;
	reg [7:0] rf_filter_coeff220_a;
	reg [7:0] rf_filter_coeff220_b;
	reg [7:0] rf_filter_coeff221_a;
	reg [7:0] rf_filter_coeff221_b;
	reg [7:0] rf_filter_coeff222_a;
	reg [7:0] rf_filter_coeff222_b;
	reg [7:0] rf_filter_coeff223_a;
	reg [7:0] rf_filter_coeff223_b;
	reg [7:0] rf_filter_coeff224_a;
	reg [7:0] rf_filter_coeff224_b;
	reg [7:0] rf_filter_coeff225_a;
	reg [7:0] rf_filter_coeff225_b;
	reg [7:0] rf_filter_coeff226_a;
	reg [7:0] rf_filter_coeff226_b;
	reg [7:0] rf_filter_coeff227_a;
	reg [7:0] rf_filter_coeff227_b;
	reg [7:0] rf_filter_coeff228_a;
	reg [7:0] rf_filter_coeff228_b;
	reg [7:0] rf_filter_coeff229_a;
	reg [7:0] rf_filter_coeff229_b;
	reg [7:0] rf_filter_coeff230_a;
	reg [7:0] rf_filter_coeff230_b;
	reg [7:0] rf_filter_coeff231_a;
	reg [7:0] rf_filter_coeff231_b;
	reg [7:0] rf_filter_coeff232_a;
	reg [7:0] rf_filter_coeff232_b;
	reg [7:0] rf_filter_coeff233_a;
	reg [7:0] rf_filter_coeff233_b;
	reg [7:0] rf_filter_coeff234_a;
	reg [7:0] rf_filter_coeff234_b;
	reg [7:0] rf_filter_coeff235_a;
	reg [7:0] rf_filter_coeff235_b;
	reg [7:0] rf_filter_coeff236_a;
	reg [7:0] rf_filter_coeff236_b;
	reg [7:0] rf_filter_coeff237_a;
	reg [7:0] rf_filter_coeff237_b;
	reg [7:0] rf_filter_coeff238_a;
	reg [7:0] rf_filter_coeff238_b;
	reg [7:0] rf_filter_coeff239_a;
	reg [7:0] rf_filter_coeff239_b;
	reg [7:0] rf_filter_coeff240_a;
	reg [7:0] rf_filter_coeff240_b;
	reg [7:0] rf_filter_coeff241_a;
	reg [7:0] rf_filter_coeff241_b;
	reg [7:0] rf_filter_coeff242_a;
	reg [7:0] rf_filter_coeff242_b;
	reg [7:0] rf_filter_coeff243_a;
	reg [7:0] rf_filter_coeff243_b;
	reg [7:0] rf_filter_coeff244_a;
	reg [7:0] rf_filter_coeff244_b;
	reg [7:0] rf_filter_coeff245_a;
	reg [7:0] rf_filter_coeff245_b;
	reg [7:0] rf_filter_coeff246_a;
	reg [7:0] rf_filter_coeff246_b;
	reg [7:0] rf_filter_coeff247_a;
	reg [7:0] rf_filter_coeff247_b;
	reg [7:0] rf_filter_coeff248_a;
	reg [7:0] rf_filter_coeff248_b;
	reg [7:0] rf_filter_coeff249_a;
	reg [7:0] rf_filter_coeff249_b;
	reg [7:0] rf_filter_coeff250_a;
	reg [7:0] rf_filter_coeff250_b;
	reg [7:0] rf_filter_coeff251_a;
	reg [7:0] rf_filter_coeff251_b;
	reg [7:0] rf_filter_coeff252_a;
	reg [7:0] rf_filter_coeff252_b;
	reg [7:0] rf_filter_coeff253_a;
	reg [7:0] rf_filter_coeff253_b;
	reg [7:0] rf_filter_coeff254_a;
	reg [7:0] rf_filter_coeff254_b;
	reg [7:0] rf_filter_coeff255_a;
	reg [7:0] rf_filter_coeff255_b;
	reg [7:0] rf_filter_coeff256_a;
	reg [7:0] rf_filter_coeff256_b;
	reg [7:0] rf_filter_coeff257_a;
	reg [7:0] rf_filter_coeff257_b;
	reg [7:0] rf_filter_coeff258_a;
	reg [7:0] rf_filter_coeff258_b;
	reg [7:0] rf_filter_coeff259_a;
	reg [7:0] rf_filter_coeff259_b;
	reg [7:0] rf_filter_coeff260_a;
	reg [7:0] rf_filter_coeff260_b;
	reg [7:0] rf_filter_coeff261_a;
	reg [7:0] rf_filter_coeff261_b;
	reg [7:0] rf_filter_coeff262_a;
	reg [7:0] rf_filter_coeff262_b;
	reg [7:0] rf_filter_coeff263_a;
	reg [7:0] rf_filter_coeff263_b;
	reg [7:0] rf_filter_coeff264_a;
	reg [7:0] rf_filter_coeff264_b;
	reg [7:0] rf_filter_coeff265_a;
	reg [7:0] rf_filter_coeff265_b;
	reg [7:0] rf_filter_coeff266_a;
	reg [7:0] rf_filter_coeff266_b;
	reg [7:0] rf_filter_coeff267_a;
	reg [7:0] rf_filter_coeff267_b;
	reg [7:0] rf_filter_coeff268_a;
	reg [7:0] rf_filter_coeff268_b;
	reg [7:0] rf_filter_coeff269_a;
	reg [7:0] rf_filter_coeff269_b;
	reg [7:0] rf_filter_coeff270_a;
	reg [7:0] rf_filter_coeff270_b;
	reg [7:0] rf_filter_coeff271_a;
	reg [7:0] rf_filter_coeff271_b;
	reg [7:0] rf_filter_coeff272_a;
	reg [7:0] rf_filter_coeff272_b;
	reg [7:0] rf_filter_coeff273_a;
	reg [7:0] rf_filter_coeff273_b;
	reg [7:0] rf_filter_coeff274_a;
	reg [7:0] rf_filter_coeff274_b;
	reg [7:0] rf_filter_coeff275_a;
	reg [7:0] rf_filter_coeff275_b;
	reg [7:0] rf_filter_coeff276_a;
	reg [7:0] rf_filter_coeff276_b;
	reg [7:0] rf_filter_coeff277_a;
	reg [7:0] rf_filter_coeff277_b;
	reg [7:0] rf_filter_coeff278_a;
	reg [7:0] rf_filter_coeff278_b;
	reg [7:0] rf_filter_coeff279_a;
	reg [7:0] rf_filter_coeff279_b;
	reg [7:0] rf_filter_coeff280_a;
	reg [7:0] rf_filter_coeff280_b;
	reg [7:0] rf_filter_coeff281_a;
	reg [7:0] rf_filter_coeff281_b;
	reg [7:0] rf_filter_coeff282_a;
	reg [7:0] rf_filter_coeff282_b;
	reg [7:0] rf_filter_coeff283_a;
	reg [7:0] rf_filter_coeff283_b;
	reg [7:0] rf_filter_coeff284_a;
	reg [7:0] rf_filter_coeff284_b;
	reg [7:0] rf_filter_coeff285_a;
	reg [7:0] rf_filter_coeff285_b;
	reg [7:0] rf_filter_coeff286_a;
	reg [7:0] rf_filter_coeff286_b;
	reg [7:0] rf_filter_coeff287_a;
	reg [7:0] rf_filter_coeff287_b;
	reg [7:0] rf_filter_coeff288_a;
	reg [7:0] rf_filter_coeff288_b;
	reg [7:0] rf_filter_coeff289_a;
	reg [7:0] rf_filter_coeff289_b;
	reg [7:0] rf_filter_coeff290_a;
	reg [7:0] rf_filter_coeff290_b;
	reg [7:0] rf_filter_coeff291_a;
	reg [7:0] rf_filter_coeff291_b;
	reg [7:0] rf_filter_coeff292_a;
	reg [7:0] rf_filter_coeff292_b;
	reg [7:0] rf_filter_coeff293_a;
	reg [7:0] rf_filter_coeff293_b;
	reg [7:0] rf_filter_coeff294_a;
	reg [7:0] rf_filter_coeff294_b;
	reg [7:0] rf_filter_coeff295_a;
	reg [7:0] rf_filter_coeff295_b;
	reg [7:0] rf_filter_coeff296_a;
	reg [7:0] rf_filter_coeff296_b;
	reg [7:0] rf_filter_coeff297_a;
	reg [7:0] rf_filter_coeff297_b;
	reg [7:0] rf_filter_coeff298_a;
	reg [7:0] rf_filter_coeff298_b;
	reg [7:0] rf_filter_coeff299_a;
	reg [7:0] rf_filter_coeff299_b;
	reg [7:0] rf_filter_coeff300_a;
	reg [7:0] rf_filter_coeff300_b;
	reg [7:0] rf_filter_coeff301_a;
	reg [7:0] rf_filter_coeff301_b;
	reg [7:0] rf_filter_coeff302_a;
	reg [7:0] rf_filter_coeff302_b;
	reg [7:0] rf_filter_coeff303_a;
	reg [7:0] rf_filter_coeff303_b;
	reg [7:0] rf_filter_coeff304_a;
	reg [7:0] rf_filter_coeff304_b;
	reg [7:0] rf_filter_coeff305_a;
	reg [7:0] rf_filter_coeff305_b;
	reg [7:0] rf_filter_coeff306_a;
	reg [7:0] rf_filter_coeff306_b;
	reg [7:0] rf_filter_coeff307_a;
	reg [7:0] rf_filter_coeff307_b;
	reg [7:0] rf_filter_coeff308_a;
	reg [7:0] rf_filter_coeff308_b;
	reg [7:0] rf_filter_coeff309_a;
	reg [7:0] rf_filter_coeff309_b;
	reg [7:0] rf_filter_coeff310_a;
	reg [7:0] rf_filter_coeff310_b;
	reg [7:0] rf_filter_coeff311_a;
	reg [7:0] rf_filter_coeff311_b;
	reg [7:0] rf_filter_coeff312_a;
	reg [7:0] rf_filter_coeff312_b;
	reg [7:0] rf_filter_coeff313_a;
	reg [7:0] rf_filter_coeff313_b;
	reg [7:0] rf_filter_coeff314_a;
	reg [7:0] rf_filter_coeff314_b;
	reg [7:0] rf_filter_coeff315_a;
	reg [7:0] rf_filter_coeff315_b;
	reg [7:0] rf_filter_coeff316_a;
	reg [7:0] rf_filter_coeff316_b;
	reg [7:0] rf_filter_coeff317_a;
	reg [7:0] rf_filter_coeff317_b;
	reg [7:0] rf_filter_coeff318_a;
	reg [7:0] rf_filter_coeff318_b;
	reg [7:0] rf_filter_coeff319_a;
	reg [7:0] rf_filter_coeff319_b;
	reg [7:0] rf_filter_coeff320_a;
	reg [7:0] rf_filter_coeff320_b;
	reg [7:0] rf_filter_coeff321_a;
	reg [7:0] rf_filter_coeff321_b;
	reg [7:0] rf_filter_coeff322_a;
	reg [7:0] rf_filter_coeff322_b;
	reg [7:0] rf_filter_coeff323_a;
	reg [7:0] rf_filter_coeff323_b;
	reg [7:0] rf_filter_coeff324_a;
	reg [7:0] rf_filter_coeff324_b;
	reg [7:0] rf_filter_coeff325_a;
	reg [7:0] rf_filter_coeff325_b;
	reg [7:0] rf_filter_coeff326_a;
	reg [7:0] rf_filter_coeff326_b;
	reg [7:0] rf_filter_coeff327_a;
	reg [7:0] rf_filter_coeff327_b;
	reg [7:0] rf_filter_coeff328_a;
	reg [7:0] rf_filter_coeff328_b;
	reg [7:0] rf_filter_coeff329_a;
	reg [7:0] rf_filter_coeff329_b;
	reg [7:0] rf_filter_coeff330_a;
	reg [7:0] rf_filter_coeff330_b;
	reg [7:0] rf_filter_coeff331_a;
	reg [7:0] rf_filter_coeff331_b;
	reg [7:0] rf_filter_coeff332_a;
	reg [7:0] rf_filter_coeff332_b;
	reg [7:0] rf_filter_coeff333_a;
	reg [7:0] rf_filter_coeff333_b;
	reg [7:0] rf_filter_coeff334_a;
	reg [7:0] rf_filter_coeff334_b;
	reg [7:0] rf_filter_coeff335_a;
	reg [7:0] rf_filter_coeff335_b;
	reg [7:0] rf_filter_coeff336_a;
	reg [7:0] rf_filter_coeff336_b;
	reg [7:0] rf_filter_coeff337_a;
	reg [7:0] rf_filter_coeff337_b;
	reg [7:0] rf_filter_coeff338_a;
	reg [7:0] rf_filter_coeff338_b;
	reg [7:0] rf_filter_coeff339_a;
	reg [7:0] rf_filter_coeff339_b;
	reg [7:0] rf_filter_coeff340_a;
	reg [7:0] rf_filter_coeff340_b;
	reg [7:0] rf_filter_coeff341_a;
	reg [7:0] rf_filter_coeff341_b;
	reg [7:0] rf_filter_coeff342_a;
	reg [7:0] rf_filter_coeff342_b;
	reg [7:0] rf_filter_coeff343_a;
	reg [7:0] rf_filter_coeff343_b;
	reg [7:0] rf_filter_coeff344_a;
	reg [7:0] rf_filter_coeff344_b;
	reg [7:0] rf_filter_coeff345_a;
	reg [7:0] rf_filter_coeff345_b;
	reg [7:0] rf_filter_coeff346_a;
	reg [7:0] rf_filter_coeff346_b;
	reg [7:0] rf_filter_coeff347_a;
	reg [7:0] rf_filter_coeff347_b;
	reg [7:0] rf_filter_coeff348_a;
	reg [7:0] rf_filter_coeff348_b;
	reg [7:0] rf_filter_coeff349_a;
	reg [7:0] rf_filter_coeff349_b;
	reg [7:0] rf_filter_coeff350_a;
	reg [7:0] rf_filter_coeff350_b;
	reg [7:0] rf_filter_coeff351_a;
	reg [7:0] rf_filter_coeff351_b;
	reg [7:0] rf_filter_coeff352_a;
	reg [7:0] rf_filter_coeff352_b;
	reg [7:0] rf_filter_coeff353_a;
	reg [7:0] rf_filter_coeff353_b;
	reg [7:0] rf_filter_coeff354_a;
	reg [7:0] rf_filter_coeff354_b;
	reg [7:0] rf_filter_coeff355_a;
	reg [7:0] rf_filter_coeff355_b;
	reg [7:0] rf_filter_coeff356_a;
	reg [7:0] rf_filter_coeff356_b;
	reg [7:0] rf_filter_coeff357_a;
	reg [7:0] rf_filter_coeff357_b;
	reg [7:0] rf_filter_coeff358_a;
	reg [7:0] rf_filter_coeff358_b;
	reg [7:0] rf_filter_coeff359_a;
	reg [7:0] rf_filter_coeff359_b;
	reg [7:0] rf_filter_coeff360_a;
	reg [7:0] rf_filter_coeff360_b;
	reg [7:0] rf_filter_coeff361_a;
	reg [7:0] rf_filter_coeff361_b;
	reg [7:0] rf_filter_coeff362_a;
	reg [7:0] rf_filter_coeff362_b;
	reg [7:0] rf_filter_coeff363_a;
	reg [7:0] rf_filter_coeff363_b;
	reg [7:0] rf_filter_coeff364_a;
	reg [7:0] rf_filter_coeff364_b;
	reg [7:0] rf_filter_coeff365_a;
	reg [7:0] rf_filter_coeff365_b;
	reg [7:0] rf_filter_coeff366_a;
	reg [7:0] rf_filter_coeff366_b;
	reg [7:0] rf_filter_coeff367_a;
	reg [7:0] rf_filter_coeff367_b;
	reg [7:0] rf_filter_coeff368_a;
	reg [7:0] rf_filter_coeff368_b;
	reg [7:0] rf_filter_coeff369_a;
	reg [7:0] rf_filter_coeff369_b;
	reg [7:0] rf_filter_coeff370_a;
	reg [7:0] rf_filter_coeff370_b;
	reg [7:0] rf_filter_coeff371_a;
	reg [7:0] rf_filter_coeff371_b;
	reg [7:0] rf_filter_coeff372_a;
	reg [7:0] rf_filter_coeff372_b;
	reg [7:0] rf_filter_coeff373_a;
	reg [7:0] rf_filter_coeff373_b;
	reg [7:0] rf_filter_coeff374_a;
	reg [7:0] rf_filter_coeff374_b;
	reg [7:0] rf_filter_coeff375_a;
	reg [7:0] rf_filter_coeff375_b;
	reg [7:0] rf_filter_coeff376_a;
	reg [7:0] rf_filter_coeff376_b;
	reg [7:0] rf_filter_coeff377_a;
	reg [7:0] rf_filter_coeff377_b;
	reg [7:0] rf_filter_coeff378_a;
	reg [7:0] rf_filter_coeff378_b;
	reg [7:0] rf_filter_coeff379_a;
	reg [7:0] rf_filter_coeff379_b;
	reg [7:0] rf_filter_coeff380_a;
	reg [7:0] rf_filter_coeff380_b;
	reg [7:0] rf_filter_coeff381_a;
	reg [7:0] rf_filter_coeff381_b;
	reg [7:0] rf_filter_coeff382_a;
	reg [7:0] rf_filter_coeff382_b;
	reg [7:0] rf_filter_coeff383_a;
	reg [7:0] rf_filter_coeff383_b;
	reg [7:0] rf_filter_coeff384_a;
	reg [7:0] rf_filter_coeff384_b;
	reg [7:0] rf_filter_coeff385_a;
	reg [7:0] rf_filter_coeff385_b;
	reg [7:0] rf_filter_coeff386_a;
	reg [7:0] rf_filter_coeff386_b;
	reg [7:0] rf_filter_coeff387_a;
	reg [7:0] rf_filter_coeff387_b;
	reg [7:0] rf_filter_coeff388_a;
	reg [7:0] rf_filter_coeff388_b;
	reg [7:0] rf_filter_coeff389_a;
	reg [7:0] rf_filter_coeff389_b;
	reg [7:0] rf_filter_coeff390_a;
	reg [7:0] rf_filter_coeff390_b;
	reg [7:0] rf_filter_coeff391_a;
	reg [7:0] rf_filter_coeff391_b;
	reg [7:0] rf_filter_coeff392_a;
	reg [7:0] rf_filter_coeff392_b;
	reg [7:0] rf_filter_coeff393_a;
	reg [7:0] rf_filter_coeff393_b;
	reg [7:0] rf_filter_coeff394_a;
	reg [7:0] rf_filter_coeff394_b;
	reg [7:0] rf_filter_coeff395_a;
	reg [7:0] rf_filter_coeff395_b;
	reg [7:0] rf_filter_coeff396_a;
	reg [7:0] rf_filter_coeff396_b;
	reg [7:0] rf_filter_coeff397_a;
	reg [7:0] rf_filter_coeff397_b;
	reg [7:0] rf_filter_coeff398_a;
	reg [7:0] rf_filter_coeff398_b;
	reg [7:0] rf_filter_coeff399_a;
	reg [7:0] rf_filter_coeff399_b;
	reg [7:0] rf_filter_coeff400_a;
	reg [7:0] rf_filter_coeff400_b;
	reg [7:0] rf_filter_coeff401_a;
	reg [7:0] rf_filter_coeff401_b;
	reg [7:0] rf_filter_coeff402_a;
	reg [7:0] rf_filter_coeff402_b;
	reg [7:0] rf_filter_coeff403_a;
	reg [7:0] rf_filter_coeff403_b;
	reg [7:0] rf_filter_coeff404_a;
	reg [7:0] rf_filter_coeff404_b;
	reg [7:0] rf_filter_coeff405_a;
	reg [7:0] rf_filter_coeff405_b;
	reg [7:0] rf_filter_coeff406_a;
	reg [7:0] rf_filter_coeff406_b;
	reg [7:0] rf_filter_coeff407_a;
	reg [7:0] rf_filter_coeff407_b;
	reg [7:0] rf_filter_coeff408_a;
	reg [7:0] rf_filter_coeff408_b;
	reg [7:0] rf_filter_coeff409_a;
	reg [7:0] rf_filter_coeff409_b;
	reg [7:0] rf_filter_coeff410_a;
	reg [7:0] rf_filter_coeff410_b;
	reg [7:0] rf_filter_coeff411_a;
	reg [7:0] rf_filter_coeff411_b;
	reg [7:0] rf_filter_coeff412_a;
	reg [7:0] rf_filter_coeff412_b;
	reg [7:0] rf_filter_coeff413_a;
	reg [7:0] rf_filter_coeff413_b;
	reg [7:0] rf_filter_coeff414_a;
	reg [7:0] rf_filter_coeff414_b;
	reg [7:0] rf_filter_coeff415_a;
	reg [7:0] rf_filter_coeff415_b;
	reg [7:0] rf_filter_coeff416_a;
	reg [7:0] rf_filter_coeff416_b;
	reg [7:0] rf_filter_coeff417_a;
	reg [7:0] rf_filter_coeff417_b;
	reg [7:0] rf_filter_coeff418_a;
	reg [7:0] rf_filter_coeff418_b;
	reg [7:0] rf_filter_coeff419_a;
	reg [7:0] rf_filter_coeff419_b;
	reg [7:0] rf_filter_coeff420_a;
	reg [7:0] rf_filter_coeff420_b;
	reg [7:0] rf_filter_coeff421_a;
	reg [7:0] rf_filter_coeff421_b;
	reg [7:0] rf_filter_coeff422_a;
	reg [7:0] rf_filter_coeff422_b;
	reg [7:0] rf_filter_coeff423_a;
	reg [7:0] rf_filter_coeff423_b;
	reg [7:0] rf_filter_coeff424_a;
	reg [7:0] rf_filter_coeff424_b;
	reg [7:0] rf_filter_coeff425_a;
	reg [7:0] rf_filter_coeff425_b;
	reg [7:0] rf_filter_coeff426_a;
	reg [7:0] rf_filter_coeff426_b;
	reg [7:0] rf_filter_coeff427_a;
	reg [7:0] rf_filter_coeff427_b;
	reg [7:0] rf_filter_coeff428_a;
	reg [7:0] rf_filter_coeff428_b;
	reg [7:0] rf_filter_coeff429_a;
	reg [7:0] rf_filter_coeff429_b;
	reg [7:0] rf_filter_coeff430_a;
	reg [7:0] rf_filter_coeff430_b;
	reg [7:0] rf_filter_coeff431_a;
	reg [7:0] rf_filter_coeff431_b;
	reg [7:0] rf_filter_coeff432_a;
	reg [7:0] rf_filter_coeff432_b;
	reg [7:0] rf_filter_coeff433_a;
	reg [7:0] rf_filter_coeff433_b;
	reg [7:0] rf_filter_coeff434_a;
	reg [7:0] rf_filter_coeff434_b;
	reg [7:0] rf_filter_coeff435_a;
	reg [7:0] rf_filter_coeff435_b;
	reg [7:0] rf_filter_coeff436_a;
	reg [7:0] rf_filter_coeff436_b;
	reg [7:0] rf_filter_coeff437_a;
	reg [7:0] rf_filter_coeff437_b;
	reg [7:0] rf_filter_coeff438_a;
	reg [7:0] rf_filter_coeff438_b;
	reg [7:0] rf_filter_coeff439_a;
	reg [7:0] rf_filter_coeff439_b;
	reg [7:0] rf_filter_coeff440_a;
	reg [7:0] rf_filter_coeff440_b;
	reg [7:0] rf_filter_coeff441_a;
	reg [7:0] rf_filter_coeff441_b;
	reg [7:0] rf_filter_coeff442_a;
	reg [7:0] rf_filter_coeff442_b;
	reg [7:0] rf_filter_coeff443_a;
	reg [7:0] rf_filter_coeff443_b;
	reg [7:0] rf_filter_coeff444_a;
	reg [7:0] rf_filter_coeff444_b;
	reg [7:0] rf_filter_coeff445_a;
	reg [7:0] rf_filter_coeff445_b;
	reg [7:0] rf_filter_coeff446_a;
	reg [7:0] rf_filter_coeff446_b;
	reg [7:0] rf_filter_coeff447_a;
	reg [7:0] rf_filter_coeff447_b;
	reg [7:0] rf_filter_coeff448_a;
	reg [7:0] rf_filter_coeff448_b;
	reg [7:0] rf_filter_coeff449_a;
	reg [7:0] rf_filter_coeff449_b;
	reg [7:0] rf_filter_coeff450_a;
	reg [7:0] rf_filter_coeff450_b;
	reg [7:0] rf_filter_coeff451_a;
	reg [7:0] rf_filter_coeff451_b;
	reg [7:0] rf_filter_coeff452_a;
	reg [7:0] rf_filter_coeff452_b;
	reg [7:0] rf_filter_coeff453_a;
	reg [7:0] rf_filter_coeff453_b;
	reg [7:0] rf_filter_coeff454_a;
	reg [7:0] rf_filter_coeff454_b;
	reg [7:0] rf_filter_coeff455_a;
	reg [7:0] rf_filter_coeff455_b;
	reg [7:0] rf_filter_coeff456_a;
	reg [7:0] rf_filter_coeff456_b;
	reg [7:0] rf_filter_coeff457_a;
	reg [7:0] rf_filter_coeff457_b;
	reg [7:0] rf_filter_coeff458_a;
	reg [7:0] rf_filter_coeff458_b;
	reg [7:0] rf_filter_coeff459_a;
	reg [7:0] rf_filter_coeff459_b;
	reg [7:0] rf_filter_coeff460_a;
	reg [7:0] rf_filter_coeff460_b;
	reg [7:0] rf_filter_coeff461_a;
	reg [7:0] rf_filter_coeff461_b;
	reg [7:0] rf_filter_coeff462_a;
	reg [7:0] rf_filter_coeff462_b;
	reg [7:0] rf_filter_coeff463_a;
	reg [7:0] rf_filter_coeff463_b;
	reg [7:0] rf_filter_coeff464_a;
	reg [7:0] rf_filter_coeff464_b;
	reg [7:0] rf_filter_coeff465_a;
	reg [7:0] rf_filter_coeff465_b;
	reg [7:0] rf_filter_coeff466_a;
	reg [7:0] rf_filter_coeff466_b;
	reg [7:0] rf_filter_coeff467_a;
	reg [7:0] rf_filter_coeff467_b;
	reg [7:0] rf_filter_coeff468_a;
	reg [7:0] rf_filter_coeff468_b;
	reg [7:0] rf_filter_coeff469_a;
	reg [7:0] rf_filter_coeff469_b;
	reg [7:0] rf_filter_coeff470_a;
	reg [7:0] rf_filter_coeff470_b;
	reg [7:0] rf_filter_coeff471_a;
	reg [7:0] rf_filter_coeff471_b;
	reg [7:0] rf_filter_coeff472_a;
	reg [7:0] rf_filter_coeff472_b;
	reg [7:0] rf_filter_coeff473_a;
	reg [7:0] rf_filter_coeff473_b;
	reg [7:0] rf_filter_coeff474_a;
	reg [7:0] rf_filter_coeff474_b;
	reg [7:0] rf_filter_coeff475_a;
	reg [7:0] rf_filter_coeff475_b;
	reg [7:0] rf_filter_coeff476_a;
	reg [7:0] rf_filter_coeff476_b;
	reg [7:0] rf_filter_coeff477_a;
	reg [7:0] rf_filter_coeff477_b;
	reg [7:0] rf_filter_coeff478_a;
	reg [7:0] rf_filter_coeff478_b;
	reg [7:0] rf_filter_coeff479_a;
	reg [7:0] rf_filter_coeff479_b;
	reg [7:0] rf_filter_coeff480_a;
	reg [7:0] rf_filter_coeff480_b;
	reg [7:0] rf_filter_coeff481_a;
	reg [7:0] rf_filter_coeff481_b;
	reg [7:0] rf_filter_coeff482_a;
	reg [7:0] rf_filter_coeff482_b;
	reg [7:0] rf_filter_coeff483_a;
	reg [7:0] rf_filter_coeff483_b;
	reg [7:0] rf_filter_coeff484_a;
	reg [7:0] rf_filter_coeff484_b;
	reg [7:0] rf_filter_coeff485_a;
	reg [7:0] rf_filter_coeff485_b;
	reg [7:0] rf_filter_coeff486_a;
	reg [7:0] rf_filter_coeff486_b;
	reg [7:0] rf_filter_coeff487_a;
	reg [7:0] rf_filter_coeff487_b;
	reg [7:0] rf_filter_coeff488_a;
	reg [7:0] rf_filter_coeff488_b;
	reg [7:0] rf_filter_coeff489_a;
	reg [7:0] rf_filter_coeff489_b;
	reg [7:0] rf_filter_coeff490_a;
	reg [7:0] rf_filter_coeff490_b;
	reg [7:0] rf_filter_coeff491_a;
	reg [7:0] rf_filter_coeff491_b;
	reg [7:0] rf_filter_coeff492_a;
	reg [7:0] rf_filter_coeff492_b;
	reg [7:0] rf_filter_coeff493_a;
	reg [7:0] rf_filter_coeff493_b;
	reg [7:0] rf_filter_coeff494_a;
	reg [7:0] rf_filter_coeff494_b;
	reg [7:0] rf_filter_coeff495_a;
	reg [7:0] rf_filter_coeff495_b;
	reg [7:0] rf_filter_coeff496_a;
	reg [7:0] rf_filter_coeff496_b;
	reg [7:0] rf_filter_coeff497_a;
	reg [7:0] rf_filter_coeff497_b;
	reg [7:0] rf_filter_coeff498_a;
	reg [7:0] rf_filter_coeff498_b;
	reg [7:0] rf_filter_coeff499_a;
	reg [7:0] rf_filter_coeff499_b;
	reg [7:0] rf_filter_coeff500_a;
	reg [7:0] rf_filter_coeff500_b;
	reg [7:0] rf_filter_coeff501_a;
	reg [7:0] rf_filter_coeff501_b;
	reg [7:0] rf_filter_coeff502_a;
	reg [7:0] rf_filter_coeff502_b;
	reg [7:0] rf_filter_coeff503_a;
	reg [7:0] rf_filter_coeff503_b;
	reg [7:0] rf_filter_coeff504_a;
	reg [7:0] rf_filter_coeff504_b;
	reg [7:0] rf_filter_coeff505_a;
	reg [7:0] rf_filter_coeff505_b;
	reg [7:0] rf_filter_coeff506_a;
	reg [7:0] rf_filter_coeff506_b;
	reg [7:0] rf_filter_coeff507_a;
	reg [7:0] rf_filter_coeff507_b;
	reg [7:0] rf_filter_coeff508_a;
	reg [7:0] rf_filter_coeff508_b;
	reg [7:0] rf_filter_coeff509_a;
	reg [7:0] rf_filter_coeff509_b;
	reg [7:0] rf_filter_coeff510_a;
	reg [7:0] rf_filter_coeff510_b;
	reg [7:0] rf_filter_coeff511_a;
	reg [7:0] rf_filter_coeff511_b;

	// Outputs
	wire aud_in_rtr;
	wire [31:0] filt_out_data;
	wire aud_out_rts;
	wire ro_filter_ovf_flag;

	// Instantiate the Unit Under Test (UUT)
	filter uut (
		.clk(clk), 
		.rstb(rstb), 
		.filt_input_data(filt_input_data), 
		.aud_in_rts(aud_in_rts), 
		.aud_in_rtr(aud_in_rtr), 
		.filt_out_data(filt_out_data), 
		.aud_out_rts(aud_out_rts), 
		.aud_out_rtr(aud_out_rtr), 
		.rf_filter_shift(rf_filter_shift), 
		.rf_filter_clip_en(rf_filter_clip_en), 
		.trig_filter_ovf_flag_clear(trig_filter_ovf_flag_clear), 
		.ro_filter_ovf_flag(ro_filter_ovf_flag), 
		.rf_filter_coeff0_a(rf_filter_coeff0_a), 
		.rf_filter_coeff0_b(rf_filter_coeff0_b), 
		.rf_filter_coeff1_a(rf_filter_coeff1_a), 
		.rf_filter_coeff1_b(rf_filter_coeff1_b), 
		.rf_filter_coeff2_a(rf_filter_coeff2_a), 
		.rf_filter_coeff2_b(rf_filter_coeff2_b), 
		.rf_filter_coeff3_a(rf_filter_coeff3_a), 
		.rf_filter_coeff3_b(rf_filter_coeff3_b), 
		.rf_filter_coeff4_a(rf_filter_coeff4_a), 
		.rf_filter_coeff4_b(rf_filter_coeff4_b), 
		.rf_filter_coeff5_a(rf_filter_coeff5_a), 
		.rf_filter_coeff5_b(rf_filter_coeff5_b), 
		.rf_filter_coeff6_a(rf_filter_coeff6_a), 
		.rf_filter_coeff6_b(rf_filter_coeff6_b), 
		.rf_filter_coeff7_a(rf_filter_coeff7_a), 
		.rf_filter_coeff7_b(rf_filter_coeff7_b), 
		.rf_filter_coeff8_a(rf_filter_coeff8_a), 
		.rf_filter_coeff8_b(rf_filter_coeff8_b), 
		.rf_filter_coeff9_a(rf_filter_coeff9_a), 
		.rf_filter_coeff9_b(rf_filter_coeff9_b), 
		.rf_filter_coeff10_a(rf_filter_coeff10_a), 
		.rf_filter_coeff10_b(rf_filter_coeff10_b), 
		.rf_filter_coeff11_a(rf_filter_coeff11_a), 
		.rf_filter_coeff11_b(rf_filter_coeff11_b), 
		.rf_filter_coeff12_a(rf_filter_coeff12_a), 
		.rf_filter_coeff12_b(rf_filter_coeff12_b), 
		.rf_filter_coeff13_a(rf_filter_coeff13_a), 
		.rf_filter_coeff13_b(rf_filter_coeff13_b), 
		.rf_filter_coeff14_a(rf_filter_coeff14_a), 
		.rf_filter_coeff14_b(rf_filter_coeff14_b), 
		.rf_filter_coeff15_a(rf_filter_coeff15_a), 
		.rf_filter_coeff15_b(rf_filter_coeff15_b), 
		.rf_filter_coeff16_a(rf_filter_coeff16_a), 
		.rf_filter_coeff16_b(rf_filter_coeff16_b), 
		.rf_filter_coeff17_a(rf_filter_coeff17_a), 
		.rf_filter_coeff17_b(rf_filter_coeff17_b), 
		.rf_filter_coeff18_a(rf_filter_coeff18_a), 
		.rf_filter_coeff18_b(rf_filter_coeff18_b), 
		.rf_filter_coeff19_a(rf_filter_coeff19_a), 
		.rf_filter_coeff19_b(rf_filter_coeff19_b), 
		.rf_filter_coeff20_a(rf_filter_coeff20_a), 
		.rf_filter_coeff20_b(rf_filter_coeff20_b), 
		.rf_filter_coeff21_a(rf_filter_coeff21_a), 
		.rf_filter_coeff21_b(rf_filter_coeff21_b), 
		.rf_filter_coeff22_a(rf_filter_coeff22_a), 
		.rf_filter_coeff22_b(rf_filter_coeff22_b), 
		.rf_filter_coeff23_a(rf_filter_coeff23_a), 
		.rf_filter_coeff23_b(rf_filter_coeff23_b), 
		.rf_filter_coeff24_a(rf_filter_coeff24_a), 
		.rf_filter_coeff24_b(rf_filter_coeff24_b), 
		.rf_filter_coeff25_a(rf_filter_coeff25_a), 
		.rf_filter_coeff25_b(rf_filter_coeff25_b), 
		.rf_filter_coeff26_a(rf_filter_coeff26_a), 
		.rf_filter_coeff26_b(rf_filter_coeff26_b), 
		.rf_filter_coeff27_a(rf_filter_coeff27_a), 
		.rf_filter_coeff27_b(rf_filter_coeff27_b), 
		.rf_filter_coeff28_a(rf_filter_coeff28_a), 
		.rf_filter_coeff28_b(rf_filter_coeff28_b), 
		.rf_filter_coeff29_a(rf_filter_coeff29_a), 
		.rf_filter_coeff29_b(rf_filter_coeff29_b), 
		.rf_filter_coeff30_a(rf_filter_coeff30_a), 
		.rf_filter_coeff30_b(rf_filter_coeff30_b), 
		.rf_filter_coeff31_a(rf_filter_coeff31_a), 
		.rf_filter_coeff31_b(rf_filter_coeff31_b), 
		.rf_filter_coeff32_a(rf_filter_coeff32_a), 
		.rf_filter_coeff32_b(rf_filter_coeff32_b), 
		.rf_filter_coeff33_a(rf_filter_coeff33_a), 
		.rf_filter_coeff33_b(rf_filter_coeff33_b), 
		.rf_filter_coeff34_a(rf_filter_coeff34_a), 
		.rf_filter_coeff34_b(rf_filter_coeff34_b), 
		.rf_filter_coeff35_a(rf_filter_coeff35_a), 
		.rf_filter_coeff35_b(rf_filter_coeff35_b), 
		.rf_filter_coeff36_a(rf_filter_coeff36_a), 
		.rf_filter_coeff36_b(rf_filter_coeff36_b), 
		.rf_filter_coeff37_a(rf_filter_coeff37_a), 
		.rf_filter_coeff37_b(rf_filter_coeff37_b), 
		.rf_filter_coeff38_a(rf_filter_coeff38_a), 
		.rf_filter_coeff38_b(rf_filter_coeff38_b), 
		.rf_filter_coeff39_a(rf_filter_coeff39_a), 
		.rf_filter_coeff39_b(rf_filter_coeff39_b), 
		.rf_filter_coeff40_a(rf_filter_coeff40_a), 
		.rf_filter_coeff40_b(rf_filter_coeff40_b), 
		.rf_filter_coeff41_a(rf_filter_coeff41_a), 
		.rf_filter_coeff41_b(rf_filter_coeff41_b), 
		.rf_filter_coeff42_a(rf_filter_coeff42_a), 
		.rf_filter_coeff42_b(rf_filter_coeff42_b), 
		.rf_filter_coeff43_a(rf_filter_coeff43_a), 
		.rf_filter_coeff43_b(rf_filter_coeff43_b), 
		.rf_filter_coeff44_a(rf_filter_coeff44_a), 
		.rf_filter_coeff44_b(rf_filter_coeff44_b), 
		.rf_filter_coeff45_a(rf_filter_coeff45_a), 
		.rf_filter_coeff45_b(rf_filter_coeff45_b), 
		.rf_filter_coeff46_a(rf_filter_coeff46_a), 
		.rf_filter_coeff46_b(rf_filter_coeff46_b), 
		.rf_filter_coeff47_a(rf_filter_coeff47_a), 
		.rf_filter_coeff47_b(rf_filter_coeff47_b), 
		.rf_filter_coeff48_a(rf_filter_coeff48_a), 
		.rf_filter_coeff48_b(rf_filter_coeff48_b), 
		.rf_filter_coeff49_a(rf_filter_coeff49_a), 
		.rf_filter_coeff49_b(rf_filter_coeff49_b), 
		.rf_filter_coeff50_a(rf_filter_coeff50_a), 
		.rf_filter_coeff50_b(rf_filter_coeff50_b), 
		.rf_filter_coeff51_a(rf_filter_coeff51_a), 
		.rf_filter_coeff51_b(rf_filter_coeff51_b), 
		.rf_filter_coeff52_a(rf_filter_coeff52_a), 
		.rf_filter_coeff52_b(rf_filter_coeff52_b), 
		.rf_filter_coeff53_a(rf_filter_coeff53_a), 
		.rf_filter_coeff53_b(rf_filter_coeff53_b), 
		.rf_filter_coeff54_a(rf_filter_coeff54_a), 
		.rf_filter_coeff54_b(rf_filter_coeff54_b), 
		.rf_filter_coeff55_a(rf_filter_coeff55_a), 
		.rf_filter_coeff55_b(rf_filter_coeff55_b), 
		.rf_filter_coeff56_a(rf_filter_coeff56_a), 
		.rf_filter_coeff56_b(rf_filter_coeff56_b), 
		.rf_filter_coeff57_a(rf_filter_coeff57_a), 
		.rf_filter_coeff57_b(rf_filter_coeff57_b), 
		.rf_filter_coeff58_a(rf_filter_coeff58_a), 
		.rf_filter_coeff58_b(rf_filter_coeff58_b), 
		.rf_filter_coeff59_a(rf_filter_coeff59_a), 
		.rf_filter_coeff59_b(rf_filter_coeff59_b), 
		.rf_filter_coeff60_a(rf_filter_coeff60_a), 
		.rf_filter_coeff60_b(rf_filter_coeff60_b), 
		.rf_filter_coeff61_a(rf_filter_coeff61_a), 
		.rf_filter_coeff61_b(rf_filter_coeff61_b), 
		.rf_filter_coeff62_a(rf_filter_coeff62_a), 
		.rf_filter_coeff62_b(rf_filter_coeff62_b), 
		.rf_filter_coeff63_a(rf_filter_coeff63_a), 
		.rf_filter_coeff63_b(rf_filter_coeff63_b), 
		.rf_filter_coeff64_a(rf_filter_coeff64_a), 
		.rf_filter_coeff64_b(rf_filter_coeff64_b), 
		.rf_filter_coeff65_a(rf_filter_coeff65_a), 
		.rf_filter_coeff65_b(rf_filter_coeff65_b), 
		.rf_filter_coeff66_a(rf_filter_coeff66_a), 
		.rf_filter_coeff66_b(rf_filter_coeff66_b), 
		.rf_filter_coeff67_a(rf_filter_coeff67_a), 
		.rf_filter_coeff67_b(rf_filter_coeff67_b), 
		.rf_filter_coeff68_a(rf_filter_coeff68_a), 
		.rf_filter_coeff68_b(rf_filter_coeff68_b), 
		.rf_filter_coeff69_a(rf_filter_coeff69_a), 
		.rf_filter_coeff69_b(rf_filter_coeff69_b), 
		.rf_filter_coeff70_a(rf_filter_coeff70_a), 
		.rf_filter_coeff70_b(rf_filter_coeff70_b), 
		.rf_filter_coeff71_a(rf_filter_coeff71_a), 
		.rf_filter_coeff71_b(rf_filter_coeff71_b), 
		.rf_filter_coeff72_a(rf_filter_coeff72_a), 
		.rf_filter_coeff72_b(rf_filter_coeff72_b), 
		.rf_filter_coeff73_a(rf_filter_coeff73_a), 
		.rf_filter_coeff73_b(rf_filter_coeff73_b), 
		.rf_filter_coeff74_a(rf_filter_coeff74_a), 
		.rf_filter_coeff74_b(rf_filter_coeff74_b), 
		.rf_filter_coeff75_a(rf_filter_coeff75_a), 
		.rf_filter_coeff75_b(rf_filter_coeff75_b), 
		.rf_filter_coeff76_a(rf_filter_coeff76_a), 
		.rf_filter_coeff76_b(rf_filter_coeff76_b), 
		.rf_filter_coeff77_a(rf_filter_coeff77_a), 
		.rf_filter_coeff77_b(rf_filter_coeff77_b), 
		.rf_filter_coeff78_a(rf_filter_coeff78_a), 
		.rf_filter_coeff78_b(rf_filter_coeff78_b), 
		.rf_filter_coeff79_a(rf_filter_coeff79_a), 
		.rf_filter_coeff79_b(rf_filter_coeff79_b), 
		.rf_filter_coeff80_a(rf_filter_coeff80_a), 
		.rf_filter_coeff80_b(rf_filter_coeff80_b), 
		.rf_filter_coeff81_a(rf_filter_coeff81_a), 
		.rf_filter_coeff81_b(rf_filter_coeff81_b), 
		.rf_filter_coeff82_a(rf_filter_coeff82_a), 
		.rf_filter_coeff82_b(rf_filter_coeff82_b), 
		.rf_filter_coeff83_a(rf_filter_coeff83_a), 
		.rf_filter_coeff83_b(rf_filter_coeff83_b), 
		.rf_filter_coeff84_a(rf_filter_coeff84_a), 
		.rf_filter_coeff84_b(rf_filter_coeff84_b), 
		.rf_filter_coeff85_a(rf_filter_coeff85_a), 
		.rf_filter_coeff85_b(rf_filter_coeff85_b), 
		.rf_filter_coeff86_a(rf_filter_coeff86_a), 
		.rf_filter_coeff86_b(rf_filter_coeff86_b), 
		.rf_filter_coeff87_a(rf_filter_coeff87_a), 
		.rf_filter_coeff87_b(rf_filter_coeff87_b), 
		.rf_filter_coeff88_a(rf_filter_coeff88_a), 
		.rf_filter_coeff88_b(rf_filter_coeff88_b), 
		.rf_filter_coeff89_a(rf_filter_coeff89_a), 
		.rf_filter_coeff89_b(rf_filter_coeff89_b), 
		.rf_filter_coeff90_a(rf_filter_coeff90_a), 
		.rf_filter_coeff90_b(rf_filter_coeff90_b), 
		.rf_filter_coeff91_a(rf_filter_coeff91_a), 
		.rf_filter_coeff91_b(rf_filter_coeff91_b), 
		.rf_filter_coeff92_a(rf_filter_coeff92_a), 
		.rf_filter_coeff92_b(rf_filter_coeff92_b), 
		.rf_filter_coeff93_a(rf_filter_coeff93_a), 
		.rf_filter_coeff93_b(rf_filter_coeff93_b), 
		.rf_filter_coeff94_a(rf_filter_coeff94_a), 
		.rf_filter_coeff94_b(rf_filter_coeff94_b), 
		.rf_filter_coeff95_a(rf_filter_coeff95_a), 
		.rf_filter_coeff95_b(rf_filter_coeff95_b), 
		.rf_filter_coeff96_a(rf_filter_coeff96_a), 
		.rf_filter_coeff96_b(rf_filter_coeff96_b), 
		.rf_filter_coeff97_a(rf_filter_coeff97_a), 
		.rf_filter_coeff97_b(rf_filter_coeff97_b), 
		.rf_filter_coeff98_a(rf_filter_coeff98_a), 
		.rf_filter_coeff98_b(rf_filter_coeff98_b), 
		.rf_filter_coeff99_a(rf_filter_coeff99_a), 
		.rf_filter_coeff99_b(rf_filter_coeff99_b), 
		.rf_filter_coeff100_a(rf_filter_coeff100_a), 
		.rf_filter_coeff100_b(rf_filter_coeff100_b), 
		.rf_filter_coeff101_a(rf_filter_coeff101_a), 
		.rf_filter_coeff101_b(rf_filter_coeff101_b), 
		.rf_filter_coeff102_a(rf_filter_coeff102_a), 
		.rf_filter_coeff102_b(rf_filter_coeff102_b), 
		.rf_filter_coeff103_a(rf_filter_coeff103_a), 
		.rf_filter_coeff103_b(rf_filter_coeff103_b), 
		.rf_filter_coeff104_a(rf_filter_coeff104_a), 
		.rf_filter_coeff104_b(rf_filter_coeff104_b), 
		.rf_filter_coeff105_a(rf_filter_coeff105_a), 
		.rf_filter_coeff105_b(rf_filter_coeff105_b), 
		.rf_filter_coeff106_a(rf_filter_coeff106_a), 
		.rf_filter_coeff106_b(rf_filter_coeff106_b), 
		.rf_filter_coeff107_a(rf_filter_coeff107_a), 
		.rf_filter_coeff107_b(rf_filter_coeff107_b), 
		.rf_filter_coeff108_a(rf_filter_coeff108_a), 
		.rf_filter_coeff108_b(rf_filter_coeff108_b), 
		.rf_filter_coeff109_a(rf_filter_coeff109_a), 
		.rf_filter_coeff109_b(rf_filter_coeff109_b), 
		.rf_filter_coeff110_a(rf_filter_coeff110_a), 
		.rf_filter_coeff110_b(rf_filter_coeff110_b), 
		.rf_filter_coeff111_a(rf_filter_coeff111_a), 
		.rf_filter_coeff111_b(rf_filter_coeff111_b), 
		.rf_filter_coeff112_a(rf_filter_coeff112_a), 
		.rf_filter_coeff112_b(rf_filter_coeff112_b), 
		.rf_filter_coeff113_a(rf_filter_coeff113_a), 
		.rf_filter_coeff113_b(rf_filter_coeff113_b), 
		.rf_filter_coeff114_a(rf_filter_coeff114_a), 
		.rf_filter_coeff114_b(rf_filter_coeff114_b), 
		.rf_filter_coeff115_a(rf_filter_coeff115_a), 
		.rf_filter_coeff115_b(rf_filter_coeff115_b), 
		.rf_filter_coeff116_a(rf_filter_coeff116_a), 
		.rf_filter_coeff116_b(rf_filter_coeff116_b), 
		.rf_filter_coeff117_a(rf_filter_coeff117_a), 
		.rf_filter_coeff117_b(rf_filter_coeff117_b), 
		.rf_filter_coeff118_a(rf_filter_coeff118_a), 
		.rf_filter_coeff118_b(rf_filter_coeff118_b), 
		.rf_filter_coeff119_a(rf_filter_coeff119_a), 
		.rf_filter_coeff119_b(rf_filter_coeff119_b), 
		.rf_filter_coeff120_a(rf_filter_coeff120_a), 
		.rf_filter_coeff120_b(rf_filter_coeff120_b), 
		.rf_filter_coeff121_a(rf_filter_coeff121_a), 
		.rf_filter_coeff121_b(rf_filter_coeff121_b), 
		.rf_filter_coeff122_a(rf_filter_coeff122_a), 
		.rf_filter_coeff122_b(rf_filter_coeff122_b), 
		.rf_filter_coeff123_a(rf_filter_coeff123_a), 
		.rf_filter_coeff123_b(rf_filter_coeff123_b), 
		.rf_filter_coeff124_a(rf_filter_coeff124_a), 
		.rf_filter_coeff124_b(rf_filter_coeff124_b), 
		.rf_filter_coeff125_a(rf_filter_coeff125_a), 
		.rf_filter_coeff125_b(rf_filter_coeff125_b), 
		.rf_filter_coeff126_a(rf_filter_coeff126_a), 
		.rf_filter_coeff126_b(rf_filter_coeff126_b), 
		.rf_filter_coeff127_a(rf_filter_coeff127_a), 
		.rf_filter_coeff127_b(rf_filter_coeff127_b), 
		.rf_filter_coeff128_a(rf_filter_coeff128_a), 
		.rf_filter_coeff128_b(rf_filter_coeff128_b), 
		.rf_filter_coeff129_a(rf_filter_coeff129_a), 
		.rf_filter_coeff129_b(rf_filter_coeff129_b), 
		.rf_filter_coeff130_a(rf_filter_coeff130_a), 
		.rf_filter_coeff130_b(rf_filter_coeff130_b), 
		.rf_filter_coeff131_a(rf_filter_coeff131_a), 
		.rf_filter_coeff131_b(rf_filter_coeff131_b), 
		.rf_filter_coeff132_a(rf_filter_coeff132_a), 
		.rf_filter_coeff132_b(rf_filter_coeff132_b), 
		.rf_filter_coeff133_a(rf_filter_coeff133_a), 
		.rf_filter_coeff133_b(rf_filter_coeff133_b), 
		.rf_filter_coeff134_a(rf_filter_coeff134_a), 
		.rf_filter_coeff134_b(rf_filter_coeff134_b), 
		.rf_filter_coeff135_a(rf_filter_coeff135_a), 
		.rf_filter_coeff135_b(rf_filter_coeff135_b), 
		.rf_filter_coeff136_a(rf_filter_coeff136_a), 
		.rf_filter_coeff136_b(rf_filter_coeff136_b), 
		.rf_filter_coeff137_a(rf_filter_coeff137_a), 
		.rf_filter_coeff137_b(rf_filter_coeff137_b), 
		.rf_filter_coeff138_a(rf_filter_coeff138_a), 
		.rf_filter_coeff138_b(rf_filter_coeff138_b), 
		.rf_filter_coeff139_a(rf_filter_coeff139_a), 
		.rf_filter_coeff139_b(rf_filter_coeff139_b), 
		.rf_filter_coeff140_a(rf_filter_coeff140_a), 
		.rf_filter_coeff140_b(rf_filter_coeff140_b), 
		.rf_filter_coeff141_a(rf_filter_coeff141_a), 
		.rf_filter_coeff141_b(rf_filter_coeff141_b), 
		.rf_filter_coeff142_a(rf_filter_coeff142_a), 
		.rf_filter_coeff142_b(rf_filter_coeff142_b), 
		.rf_filter_coeff143_a(rf_filter_coeff143_a), 
		.rf_filter_coeff143_b(rf_filter_coeff143_b), 
		.rf_filter_coeff144_a(rf_filter_coeff144_a), 
		.rf_filter_coeff144_b(rf_filter_coeff144_b), 
		.rf_filter_coeff145_a(rf_filter_coeff145_a), 
		.rf_filter_coeff145_b(rf_filter_coeff145_b), 
		.rf_filter_coeff146_a(rf_filter_coeff146_a), 
		.rf_filter_coeff146_b(rf_filter_coeff146_b), 
		.rf_filter_coeff147_a(rf_filter_coeff147_a), 
		.rf_filter_coeff147_b(rf_filter_coeff147_b), 
		.rf_filter_coeff148_a(rf_filter_coeff148_a), 
		.rf_filter_coeff148_b(rf_filter_coeff148_b), 
		.rf_filter_coeff149_a(rf_filter_coeff149_a), 
		.rf_filter_coeff149_b(rf_filter_coeff149_b), 
		.rf_filter_coeff150_a(rf_filter_coeff150_a), 
		.rf_filter_coeff150_b(rf_filter_coeff150_b), 
		.rf_filter_coeff151_a(rf_filter_coeff151_a), 
		.rf_filter_coeff151_b(rf_filter_coeff151_b), 
		.rf_filter_coeff152_a(rf_filter_coeff152_a), 
		.rf_filter_coeff152_b(rf_filter_coeff152_b), 
		.rf_filter_coeff153_a(rf_filter_coeff153_a), 
		.rf_filter_coeff153_b(rf_filter_coeff153_b), 
		.rf_filter_coeff154_a(rf_filter_coeff154_a), 
		.rf_filter_coeff154_b(rf_filter_coeff154_b), 
		.rf_filter_coeff155_a(rf_filter_coeff155_a), 
		.rf_filter_coeff155_b(rf_filter_coeff155_b), 
		.rf_filter_coeff156_a(rf_filter_coeff156_a), 
		.rf_filter_coeff156_b(rf_filter_coeff156_b), 
		.rf_filter_coeff157_a(rf_filter_coeff157_a), 
		.rf_filter_coeff157_b(rf_filter_coeff157_b), 
		.rf_filter_coeff158_a(rf_filter_coeff158_a), 
		.rf_filter_coeff158_b(rf_filter_coeff158_b), 
		.rf_filter_coeff159_a(rf_filter_coeff159_a), 
		.rf_filter_coeff159_b(rf_filter_coeff159_b), 
		.rf_filter_coeff160_a(rf_filter_coeff160_a), 
		.rf_filter_coeff160_b(rf_filter_coeff160_b), 
		.rf_filter_coeff161_a(rf_filter_coeff161_a), 
		.rf_filter_coeff161_b(rf_filter_coeff161_b), 
		.rf_filter_coeff162_a(rf_filter_coeff162_a), 
		.rf_filter_coeff162_b(rf_filter_coeff162_b), 
		.rf_filter_coeff163_a(rf_filter_coeff163_a), 
		.rf_filter_coeff163_b(rf_filter_coeff163_b), 
		.rf_filter_coeff164_a(rf_filter_coeff164_a), 
		.rf_filter_coeff164_b(rf_filter_coeff164_b), 
		.rf_filter_coeff165_a(rf_filter_coeff165_a), 
		.rf_filter_coeff165_b(rf_filter_coeff165_b), 
		.rf_filter_coeff166_a(rf_filter_coeff166_a), 
		.rf_filter_coeff166_b(rf_filter_coeff166_b), 
		.rf_filter_coeff167_a(rf_filter_coeff167_a), 
		.rf_filter_coeff167_b(rf_filter_coeff167_b), 
		.rf_filter_coeff168_a(rf_filter_coeff168_a), 
		.rf_filter_coeff168_b(rf_filter_coeff168_b), 
		.rf_filter_coeff169_a(rf_filter_coeff169_a), 
		.rf_filter_coeff169_b(rf_filter_coeff169_b), 
		.rf_filter_coeff170_a(rf_filter_coeff170_a), 
		.rf_filter_coeff170_b(rf_filter_coeff170_b), 
		.rf_filter_coeff171_a(rf_filter_coeff171_a), 
		.rf_filter_coeff171_b(rf_filter_coeff171_b), 
		.rf_filter_coeff172_a(rf_filter_coeff172_a), 
		.rf_filter_coeff172_b(rf_filter_coeff172_b), 
		.rf_filter_coeff173_a(rf_filter_coeff173_a), 
		.rf_filter_coeff173_b(rf_filter_coeff173_b), 
		.rf_filter_coeff174_a(rf_filter_coeff174_a), 
		.rf_filter_coeff174_b(rf_filter_coeff174_b), 
		.rf_filter_coeff175_a(rf_filter_coeff175_a), 
		.rf_filter_coeff175_b(rf_filter_coeff175_b), 
		.rf_filter_coeff176_a(rf_filter_coeff176_a), 
		.rf_filter_coeff176_b(rf_filter_coeff176_b), 
		.rf_filter_coeff177_a(rf_filter_coeff177_a), 
		.rf_filter_coeff177_b(rf_filter_coeff177_b), 
		.rf_filter_coeff178_a(rf_filter_coeff178_a), 
		.rf_filter_coeff178_b(rf_filter_coeff178_b), 
		.rf_filter_coeff179_a(rf_filter_coeff179_a), 
		.rf_filter_coeff179_b(rf_filter_coeff179_b), 
		.rf_filter_coeff180_a(rf_filter_coeff180_a), 
		.rf_filter_coeff180_b(rf_filter_coeff180_b), 
		.rf_filter_coeff181_a(rf_filter_coeff181_a), 
		.rf_filter_coeff181_b(rf_filter_coeff181_b), 
		.rf_filter_coeff182_a(rf_filter_coeff182_a), 
		.rf_filter_coeff182_b(rf_filter_coeff182_b), 
		.rf_filter_coeff183_a(rf_filter_coeff183_a), 
		.rf_filter_coeff183_b(rf_filter_coeff183_b), 
		.rf_filter_coeff184_a(rf_filter_coeff184_a), 
		.rf_filter_coeff184_b(rf_filter_coeff184_b), 
		.rf_filter_coeff185_a(rf_filter_coeff185_a), 
		.rf_filter_coeff185_b(rf_filter_coeff185_b), 
		.rf_filter_coeff186_a(rf_filter_coeff186_a), 
		.rf_filter_coeff186_b(rf_filter_coeff186_b), 
		.rf_filter_coeff187_a(rf_filter_coeff187_a), 
		.rf_filter_coeff187_b(rf_filter_coeff187_b), 
		.rf_filter_coeff188_a(rf_filter_coeff188_a), 
		.rf_filter_coeff188_b(rf_filter_coeff188_b), 
		.rf_filter_coeff189_a(rf_filter_coeff189_a), 
		.rf_filter_coeff189_b(rf_filter_coeff189_b), 
		.rf_filter_coeff190_a(rf_filter_coeff190_a), 
		.rf_filter_coeff190_b(rf_filter_coeff190_b), 
		.rf_filter_coeff191_a(rf_filter_coeff191_a), 
		.rf_filter_coeff191_b(rf_filter_coeff191_b), 
		.rf_filter_coeff192_a(rf_filter_coeff192_a), 
		.rf_filter_coeff192_b(rf_filter_coeff192_b), 
		.rf_filter_coeff193_a(rf_filter_coeff193_a), 
		.rf_filter_coeff193_b(rf_filter_coeff193_b), 
		.rf_filter_coeff194_a(rf_filter_coeff194_a), 
		.rf_filter_coeff194_b(rf_filter_coeff194_b), 
		.rf_filter_coeff195_a(rf_filter_coeff195_a), 
		.rf_filter_coeff195_b(rf_filter_coeff195_b), 
		.rf_filter_coeff196_a(rf_filter_coeff196_a), 
		.rf_filter_coeff196_b(rf_filter_coeff196_b), 
		.rf_filter_coeff197_a(rf_filter_coeff197_a), 
		.rf_filter_coeff197_b(rf_filter_coeff197_b), 
		.rf_filter_coeff198_a(rf_filter_coeff198_a), 
		.rf_filter_coeff198_b(rf_filter_coeff198_b), 
		.rf_filter_coeff199_a(rf_filter_coeff199_a), 
		.rf_filter_coeff199_b(rf_filter_coeff199_b), 
		.rf_filter_coeff200_a(rf_filter_coeff200_a), 
		.rf_filter_coeff200_b(rf_filter_coeff200_b), 
		.rf_filter_coeff201_a(rf_filter_coeff201_a), 
		.rf_filter_coeff201_b(rf_filter_coeff201_b), 
		.rf_filter_coeff202_a(rf_filter_coeff202_a), 
		.rf_filter_coeff202_b(rf_filter_coeff202_b), 
		.rf_filter_coeff203_a(rf_filter_coeff203_a), 
		.rf_filter_coeff203_b(rf_filter_coeff203_b), 
		.rf_filter_coeff204_a(rf_filter_coeff204_a), 
		.rf_filter_coeff204_b(rf_filter_coeff204_b), 
		.rf_filter_coeff205_a(rf_filter_coeff205_a), 
		.rf_filter_coeff205_b(rf_filter_coeff205_b), 
		.rf_filter_coeff206_a(rf_filter_coeff206_a), 
		.rf_filter_coeff206_b(rf_filter_coeff206_b), 
		.rf_filter_coeff207_a(rf_filter_coeff207_a), 
		.rf_filter_coeff207_b(rf_filter_coeff207_b), 
		.rf_filter_coeff208_a(rf_filter_coeff208_a), 
		.rf_filter_coeff208_b(rf_filter_coeff208_b), 
		.rf_filter_coeff209_a(rf_filter_coeff209_a), 
		.rf_filter_coeff209_b(rf_filter_coeff209_b), 
		.rf_filter_coeff210_a(rf_filter_coeff210_a), 
		.rf_filter_coeff210_b(rf_filter_coeff210_b), 
		.rf_filter_coeff211_a(rf_filter_coeff211_a), 
		.rf_filter_coeff211_b(rf_filter_coeff211_b), 
		.rf_filter_coeff212_a(rf_filter_coeff212_a), 
		.rf_filter_coeff212_b(rf_filter_coeff212_b), 
		.rf_filter_coeff213_a(rf_filter_coeff213_a), 
		.rf_filter_coeff213_b(rf_filter_coeff213_b), 
		.rf_filter_coeff214_a(rf_filter_coeff214_a), 
		.rf_filter_coeff214_b(rf_filter_coeff214_b), 
		.rf_filter_coeff215_a(rf_filter_coeff215_a), 
		.rf_filter_coeff215_b(rf_filter_coeff215_b), 
		.rf_filter_coeff216_a(rf_filter_coeff216_a), 
		.rf_filter_coeff216_b(rf_filter_coeff216_b), 
		.rf_filter_coeff217_a(rf_filter_coeff217_a), 
		.rf_filter_coeff217_b(rf_filter_coeff217_b), 
		.rf_filter_coeff218_a(rf_filter_coeff218_a), 
		.rf_filter_coeff218_b(rf_filter_coeff218_b), 
		.rf_filter_coeff219_a(rf_filter_coeff219_a), 
		.rf_filter_coeff219_b(rf_filter_coeff219_b), 
		.rf_filter_coeff220_a(rf_filter_coeff220_a), 
		.rf_filter_coeff220_b(rf_filter_coeff220_b), 
		.rf_filter_coeff221_a(rf_filter_coeff221_a), 
		.rf_filter_coeff221_b(rf_filter_coeff221_b), 
		.rf_filter_coeff222_a(rf_filter_coeff222_a), 
		.rf_filter_coeff222_b(rf_filter_coeff222_b), 
		.rf_filter_coeff223_a(rf_filter_coeff223_a), 
		.rf_filter_coeff223_b(rf_filter_coeff223_b), 
		.rf_filter_coeff224_a(rf_filter_coeff224_a), 
		.rf_filter_coeff224_b(rf_filter_coeff224_b), 
		.rf_filter_coeff225_a(rf_filter_coeff225_a), 
		.rf_filter_coeff225_b(rf_filter_coeff225_b), 
		.rf_filter_coeff226_a(rf_filter_coeff226_a), 
		.rf_filter_coeff226_b(rf_filter_coeff226_b), 
		.rf_filter_coeff227_a(rf_filter_coeff227_a), 
		.rf_filter_coeff227_b(rf_filter_coeff227_b), 
		.rf_filter_coeff228_a(rf_filter_coeff228_a), 
		.rf_filter_coeff228_b(rf_filter_coeff228_b), 
		.rf_filter_coeff229_a(rf_filter_coeff229_a), 
		.rf_filter_coeff229_b(rf_filter_coeff229_b), 
		.rf_filter_coeff230_a(rf_filter_coeff230_a), 
		.rf_filter_coeff230_b(rf_filter_coeff230_b), 
		.rf_filter_coeff231_a(rf_filter_coeff231_a), 
		.rf_filter_coeff231_b(rf_filter_coeff231_b), 
		.rf_filter_coeff232_a(rf_filter_coeff232_a), 
		.rf_filter_coeff232_b(rf_filter_coeff232_b), 
		.rf_filter_coeff233_a(rf_filter_coeff233_a), 
		.rf_filter_coeff233_b(rf_filter_coeff233_b), 
		.rf_filter_coeff234_a(rf_filter_coeff234_a), 
		.rf_filter_coeff234_b(rf_filter_coeff234_b), 
		.rf_filter_coeff235_a(rf_filter_coeff235_a), 
		.rf_filter_coeff235_b(rf_filter_coeff235_b), 
		.rf_filter_coeff236_a(rf_filter_coeff236_a), 
		.rf_filter_coeff236_b(rf_filter_coeff236_b), 
		.rf_filter_coeff237_a(rf_filter_coeff237_a), 
		.rf_filter_coeff237_b(rf_filter_coeff237_b), 
		.rf_filter_coeff238_a(rf_filter_coeff238_a), 
		.rf_filter_coeff238_b(rf_filter_coeff238_b), 
		.rf_filter_coeff239_a(rf_filter_coeff239_a), 
		.rf_filter_coeff239_b(rf_filter_coeff239_b), 
		.rf_filter_coeff240_a(rf_filter_coeff240_a), 
		.rf_filter_coeff240_b(rf_filter_coeff240_b), 
		.rf_filter_coeff241_a(rf_filter_coeff241_a), 
		.rf_filter_coeff241_b(rf_filter_coeff241_b), 
		.rf_filter_coeff242_a(rf_filter_coeff242_a), 
		.rf_filter_coeff242_b(rf_filter_coeff242_b), 
		.rf_filter_coeff243_a(rf_filter_coeff243_a), 
		.rf_filter_coeff243_b(rf_filter_coeff243_b), 
		.rf_filter_coeff244_a(rf_filter_coeff244_a), 
		.rf_filter_coeff244_b(rf_filter_coeff244_b), 
		.rf_filter_coeff245_a(rf_filter_coeff245_a), 
		.rf_filter_coeff245_b(rf_filter_coeff245_b), 
		.rf_filter_coeff246_a(rf_filter_coeff246_a), 
		.rf_filter_coeff246_b(rf_filter_coeff246_b), 
		.rf_filter_coeff247_a(rf_filter_coeff247_a), 
		.rf_filter_coeff247_b(rf_filter_coeff247_b), 
		.rf_filter_coeff248_a(rf_filter_coeff248_a), 
		.rf_filter_coeff248_b(rf_filter_coeff248_b), 
		.rf_filter_coeff249_a(rf_filter_coeff249_a), 
		.rf_filter_coeff249_b(rf_filter_coeff249_b), 
		.rf_filter_coeff250_a(rf_filter_coeff250_a), 
		.rf_filter_coeff250_b(rf_filter_coeff250_b), 
		.rf_filter_coeff251_a(rf_filter_coeff251_a), 
		.rf_filter_coeff251_b(rf_filter_coeff251_b), 
		.rf_filter_coeff252_a(rf_filter_coeff252_a), 
		.rf_filter_coeff252_b(rf_filter_coeff252_b), 
		.rf_filter_coeff253_a(rf_filter_coeff253_a), 
		.rf_filter_coeff253_b(rf_filter_coeff253_b), 
		.rf_filter_coeff254_a(rf_filter_coeff254_a), 
		.rf_filter_coeff254_b(rf_filter_coeff254_b), 
		.rf_filter_coeff255_a(rf_filter_coeff255_a), 
		.rf_filter_coeff255_b(rf_filter_coeff255_b), 
		.rf_filter_coeff256_a(rf_filter_coeff256_a), 
		.rf_filter_coeff256_b(rf_filter_coeff256_b), 
		.rf_filter_coeff257_a(rf_filter_coeff257_a), 
		.rf_filter_coeff257_b(rf_filter_coeff257_b), 
		.rf_filter_coeff258_a(rf_filter_coeff258_a), 
		.rf_filter_coeff258_b(rf_filter_coeff258_b), 
		.rf_filter_coeff259_a(rf_filter_coeff259_a), 
		.rf_filter_coeff259_b(rf_filter_coeff259_b), 
		.rf_filter_coeff260_a(rf_filter_coeff260_a), 
		.rf_filter_coeff260_b(rf_filter_coeff260_b), 
		.rf_filter_coeff261_a(rf_filter_coeff261_a), 
		.rf_filter_coeff261_b(rf_filter_coeff261_b), 
		.rf_filter_coeff262_a(rf_filter_coeff262_a), 
		.rf_filter_coeff262_b(rf_filter_coeff262_b), 
		.rf_filter_coeff263_a(rf_filter_coeff263_a), 
		.rf_filter_coeff263_b(rf_filter_coeff263_b), 
		.rf_filter_coeff264_a(rf_filter_coeff264_a), 
		.rf_filter_coeff264_b(rf_filter_coeff264_b), 
		.rf_filter_coeff265_a(rf_filter_coeff265_a), 
		.rf_filter_coeff265_b(rf_filter_coeff265_b), 
		.rf_filter_coeff266_a(rf_filter_coeff266_a), 
		.rf_filter_coeff266_b(rf_filter_coeff266_b), 
		.rf_filter_coeff267_a(rf_filter_coeff267_a), 
		.rf_filter_coeff267_b(rf_filter_coeff267_b), 
		.rf_filter_coeff268_a(rf_filter_coeff268_a), 
		.rf_filter_coeff268_b(rf_filter_coeff268_b), 
		.rf_filter_coeff269_a(rf_filter_coeff269_a), 
		.rf_filter_coeff269_b(rf_filter_coeff269_b), 
		.rf_filter_coeff270_a(rf_filter_coeff270_a), 
		.rf_filter_coeff270_b(rf_filter_coeff270_b), 
		.rf_filter_coeff271_a(rf_filter_coeff271_a), 
		.rf_filter_coeff271_b(rf_filter_coeff271_b), 
		.rf_filter_coeff272_a(rf_filter_coeff272_a), 
		.rf_filter_coeff272_b(rf_filter_coeff272_b), 
		.rf_filter_coeff273_a(rf_filter_coeff273_a), 
		.rf_filter_coeff273_b(rf_filter_coeff273_b), 
		.rf_filter_coeff274_a(rf_filter_coeff274_a), 
		.rf_filter_coeff274_b(rf_filter_coeff274_b), 
		.rf_filter_coeff275_a(rf_filter_coeff275_a), 
		.rf_filter_coeff275_b(rf_filter_coeff275_b), 
		.rf_filter_coeff276_a(rf_filter_coeff276_a), 
		.rf_filter_coeff276_b(rf_filter_coeff276_b), 
		.rf_filter_coeff277_a(rf_filter_coeff277_a), 
		.rf_filter_coeff277_b(rf_filter_coeff277_b), 
		.rf_filter_coeff278_a(rf_filter_coeff278_a), 
		.rf_filter_coeff278_b(rf_filter_coeff278_b), 
		.rf_filter_coeff279_a(rf_filter_coeff279_a), 
		.rf_filter_coeff279_b(rf_filter_coeff279_b), 
		.rf_filter_coeff280_a(rf_filter_coeff280_a), 
		.rf_filter_coeff280_b(rf_filter_coeff280_b), 
		.rf_filter_coeff281_a(rf_filter_coeff281_a), 
		.rf_filter_coeff281_b(rf_filter_coeff281_b), 
		.rf_filter_coeff282_a(rf_filter_coeff282_a), 
		.rf_filter_coeff282_b(rf_filter_coeff282_b), 
		.rf_filter_coeff283_a(rf_filter_coeff283_a), 
		.rf_filter_coeff283_b(rf_filter_coeff283_b), 
		.rf_filter_coeff284_a(rf_filter_coeff284_a), 
		.rf_filter_coeff284_b(rf_filter_coeff284_b), 
		.rf_filter_coeff285_a(rf_filter_coeff285_a), 
		.rf_filter_coeff285_b(rf_filter_coeff285_b), 
		.rf_filter_coeff286_a(rf_filter_coeff286_a), 
		.rf_filter_coeff286_b(rf_filter_coeff286_b), 
		.rf_filter_coeff287_a(rf_filter_coeff287_a), 
		.rf_filter_coeff287_b(rf_filter_coeff287_b), 
		.rf_filter_coeff288_a(rf_filter_coeff288_a), 
		.rf_filter_coeff288_b(rf_filter_coeff288_b), 
		.rf_filter_coeff289_a(rf_filter_coeff289_a), 
		.rf_filter_coeff289_b(rf_filter_coeff289_b), 
		.rf_filter_coeff290_a(rf_filter_coeff290_a), 
		.rf_filter_coeff290_b(rf_filter_coeff290_b), 
		.rf_filter_coeff291_a(rf_filter_coeff291_a), 
		.rf_filter_coeff291_b(rf_filter_coeff291_b), 
		.rf_filter_coeff292_a(rf_filter_coeff292_a), 
		.rf_filter_coeff292_b(rf_filter_coeff292_b), 
		.rf_filter_coeff293_a(rf_filter_coeff293_a), 
		.rf_filter_coeff293_b(rf_filter_coeff293_b), 
		.rf_filter_coeff294_a(rf_filter_coeff294_a), 
		.rf_filter_coeff294_b(rf_filter_coeff294_b), 
		.rf_filter_coeff295_a(rf_filter_coeff295_a), 
		.rf_filter_coeff295_b(rf_filter_coeff295_b), 
		.rf_filter_coeff296_a(rf_filter_coeff296_a), 
		.rf_filter_coeff296_b(rf_filter_coeff296_b), 
		.rf_filter_coeff297_a(rf_filter_coeff297_a), 
		.rf_filter_coeff297_b(rf_filter_coeff297_b), 
		.rf_filter_coeff298_a(rf_filter_coeff298_a), 
		.rf_filter_coeff298_b(rf_filter_coeff298_b), 
		.rf_filter_coeff299_a(rf_filter_coeff299_a), 
		.rf_filter_coeff299_b(rf_filter_coeff299_b), 
		.rf_filter_coeff300_a(rf_filter_coeff300_a), 
		.rf_filter_coeff300_b(rf_filter_coeff300_b), 
		.rf_filter_coeff301_a(rf_filter_coeff301_a), 
		.rf_filter_coeff301_b(rf_filter_coeff301_b), 
		.rf_filter_coeff302_a(rf_filter_coeff302_a), 
		.rf_filter_coeff302_b(rf_filter_coeff302_b), 
		.rf_filter_coeff303_a(rf_filter_coeff303_a), 
		.rf_filter_coeff303_b(rf_filter_coeff303_b), 
		.rf_filter_coeff304_a(rf_filter_coeff304_a), 
		.rf_filter_coeff304_b(rf_filter_coeff304_b), 
		.rf_filter_coeff305_a(rf_filter_coeff305_a), 
		.rf_filter_coeff305_b(rf_filter_coeff305_b), 
		.rf_filter_coeff306_a(rf_filter_coeff306_a), 
		.rf_filter_coeff306_b(rf_filter_coeff306_b), 
		.rf_filter_coeff307_a(rf_filter_coeff307_a), 
		.rf_filter_coeff307_b(rf_filter_coeff307_b), 
		.rf_filter_coeff308_a(rf_filter_coeff308_a), 
		.rf_filter_coeff308_b(rf_filter_coeff308_b), 
		.rf_filter_coeff309_a(rf_filter_coeff309_a), 
		.rf_filter_coeff309_b(rf_filter_coeff309_b), 
		.rf_filter_coeff310_a(rf_filter_coeff310_a), 
		.rf_filter_coeff310_b(rf_filter_coeff310_b), 
		.rf_filter_coeff311_a(rf_filter_coeff311_a), 
		.rf_filter_coeff311_b(rf_filter_coeff311_b), 
		.rf_filter_coeff312_a(rf_filter_coeff312_a), 
		.rf_filter_coeff312_b(rf_filter_coeff312_b), 
		.rf_filter_coeff313_a(rf_filter_coeff313_a), 
		.rf_filter_coeff313_b(rf_filter_coeff313_b), 
		.rf_filter_coeff314_a(rf_filter_coeff314_a), 
		.rf_filter_coeff314_b(rf_filter_coeff314_b), 
		.rf_filter_coeff315_a(rf_filter_coeff315_a), 
		.rf_filter_coeff315_b(rf_filter_coeff315_b), 
		.rf_filter_coeff316_a(rf_filter_coeff316_a), 
		.rf_filter_coeff316_b(rf_filter_coeff316_b), 
		.rf_filter_coeff317_a(rf_filter_coeff317_a), 
		.rf_filter_coeff317_b(rf_filter_coeff317_b), 
		.rf_filter_coeff318_a(rf_filter_coeff318_a), 
		.rf_filter_coeff318_b(rf_filter_coeff318_b), 
		.rf_filter_coeff319_a(rf_filter_coeff319_a), 
		.rf_filter_coeff319_b(rf_filter_coeff319_b), 
		.rf_filter_coeff320_a(rf_filter_coeff320_a), 
		.rf_filter_coeff320_b(rf_filter_coeff320_b), 
		.rf_filter_coeff321_a(rf_filter_coeff321_a), 
		.rf_filter_coeff321_b(rf_filter_coeff321_b), 
		.rf_filter_coeff322_a(rf_filter_coeff322_a), 
		.rf_filter_coeff322_b(rf_filter_coeff322_b), 
		.rf_filter_coeff323_a(rf_filter_coeff323_a), 
		.rf_filter_coeff323_b(rf_filter_coeff323_b), 
		.rf_filter_coeff324_a(rf_filter_coeff324_a), 
		.rf_filter_coeff324_b(rf_filter_coeff324_b), 
		.rf_filter_coeff325_a(rf_filter_coeff325_a), 
		.rf_filter_coeff325_b(rf_filter_coeff325_b), 
		.rf_filter_coeff326_a(rf_filter_coeff326_a), 
		.rf_filter_coeff326_b(rf_filter_coeff326_b), 
		.rf_filter_coeff327_a(rf_filter_coeff327_a), 
		.rf_filter_coeff327_b(rf_filter_coeff327_b), 
		.rf_filter_coeff328_a(rf_filter_coeff328_a), 
		.rf_filter_coeff328_b(rf_filter_coeff328_b), 
		.rf_filter_coeff329_a(rf_filter_coeff329_a), 
		.rf_filter_coeff329_b(rf_filter_coeff329_b), 
		.rf_filter_coeff330_a(rf_filter_coeff330_a), 
		.rf_filter_coeff330_b(rf_filter_coeff330_b), 
		.rf_filter_coeff331_a(rf_filter_coeff331_a), 
		.rf_filter_coeff331_b(rf_filter_coeff331_b), 
		.rf_filter_coeff332_a(rf_filter_coeff332_a), 
		.rf_filter_coeff332_b(rf_filter_coeff332_b), 
		.rf_filter_coeff333_a(rf_filter_coeff333_a), 
		.rf_filter_coeff333_b(rf_filter_coeff333_b), 
		.rf_filter_coeff334_a(rf_filter_coeff334_a), 
		.rf_filter_coeff334_b(rf_filter_coeff334_b), 
		.rf_filter_coeff335_a(rf_filter_coeff335_a), 
		.rf_filter_coeff335_b(rf_filter_coeff335_b), 
		.rf_filter_coeff336_a(rf_filter_coeff336_a), 
		.rf_filter_coeff336_b(rf_filter_coeff336_b), 
		.rf_filter_coeff337_a(rf_filter_coeff337_a), 
		.rf_filter_coeff337_b(rf_filter_coeff337_b), 
		.rf_filter_coeff338_a(rf_filter_coeff338_a), 
		.rf_filter_coeff338_b(rf_filter_coeff338_b), 
		.rf_filter_coeff339_a(rf_filter_coeff339_a), 
		.rf_filter_coeff339_b(rf_filter_coeff339_b), 
		.rf_filter_coeff340_a(rf_filter_coeff340_a), 
		.rf_filter_coeff340_b(rf_filter_coeff340_b), 
		.rf_filter_coeff341_a(rf_filter_coeff341_a), 
		.rf_filter_coeff341_b(rf_filter_coeff341_b), 
		.rf_filter_coeff342_a(rf_filter_coeff342_a), 
		.rf_filter_coeff342_b(rf_filter_coeff342_b), 
		.rf_filter_coeff343_a(rf_filter_coeff343_a), 
		.rf_filter_coeff343_b(rf_filter_coeff343_b), 
		.rf_filter_coeff344_a(rf_filter_coeff344_a), 
		.rf_filter_coeff344_b(rf_filter_coeff344_b), 
		.rf_filter_coeff345_a(rf_filter_coeff345_a), 
		.rf_filter_coeff345_b(rf_filter_coeff345_b), 
		.rf_filter_coeff346_a(rf_filter_coeff346_a), 
		.rf_filter_coeff346_b(rf_filter_coeff346_b), 
		.rf_filter_coeff347_a(rf_filter_coeff347_a), 
		.rf_filter_coeff347_b(rf_filter_coeff347_b), 
		.rf_filter_coeff348_a(rf_filter_coeff348_a), 
		.rf_filter_coeff348_b(rf_filter_coeff348_b), 
		.rf_filter_coeff349_a(rf_filter_coeff349_a), 
		.rf_filter_coeff349_b(rf_filter_coeff349_b), 
		.rf_filter_coeff350_a(rf_filter_coeff350_a), 
		.rf_filter_coeff350_b(rf_filter_coeff350_b), 
		.rf_filter_coeff351_a(rf_filter_coeff351_a), 
		.rf_filter_coeff351_b(rf_filter_coeff351_b), 
		.rf_filter_coeff352_a(rf_filter_coeff352_a), 
		.rf_filter_coeff352_b(rf_filter_coeff352_b), 
		.rf_filter_coeff353_a(rf_filter_coeff353_a), 
		.rf_filter_coeff353_b(rf_filter_coeff353_b), 
		.rf_filter_coeff354_a(rf_filter_coeff354_a), 
		.rf_filter_coeff354_b(rf_filter_coeff354_b), 
		.rf_filter_coeff355_a(rf_filter_coeff355_a), 
		.rf_filter_coeff355_b(rf_filter_coeff355_b), 
		.rf_filter_coeff356_a(rf_filter_coeff356_a), 
		.rf_filter_coeff356_b(rf_filter_coeff356_b), 
		.rf_filter_coeff357_a(rf_filter_coeff357_a), 
		.rf_filter_coeff357_b(rf_filter_coeff357_b), 
		.rf_filter_coeff358_a(rf_filter_coeff358_a), 
		.rf_filter_coeff358_b(rf_filter_coeff358_b), 
		.rf_filter_coeff359_a(rf_filter_coeff359_a), 
		.rf_filter_coeff359_b(rf_filter_coeff359_b), 
		.rf_filter_coeff360_a(rf_filter_coeff360_a), 
		.rf_filter_coeff360_b(rf_filter_coeff360_b), 
		.rf_filter_coeff361_a(rf_filter_coeff361_a), 
		.rf_filter_coeff361_b(rf_filter_coeff361_b), 
		.rf_filter_coeff362_a(rf_filter_coeff362_a), 
		.rf_filter_coeff362_b(rf_filter_coeff362_b), 
		.rf_filter_coeff363_a(rf_filter_coeff363_a), 
		.rf_filter_coeff363_b(rf_filter_coeff363_b), 
		.rf_filter_coeff364_a(rf_filter_coeff364_a), 
		.rf_filter_coeff364_b(rf_filter_coeff364_b), 
		.rf_filter_coeff365_a(rf_filter_coeff365_a), 
		.rf_filter_coeff365_b(rf_filter_coeff365_b), 
		.rf_filter_coeff366_a(rf_filter_coeff366_a), 
		.rf_filter_coeff366_b(rf_filter_coeff366_b), 
		.rf_filter_coeff367_a(rf_filter_coeff367_a), 
		.rf_filter_coeff367_b(rf_filter_coeff367_b), 
		.rf_filter_coeff368_a(rf_filter_coeff368_a), 
		.rf_filter_coeff368_b(rf_filter_coeff368_b), 
		.rf_filter_coeff369_a(rf_filter_coeff369_a), 
		.rf_filter_coeff369_b(rf_filter_coeff369_b), 
		.rf_filter_coeff370_a(rf_filter_coeff370_a), 
		.rf_filter_coeff370_b(rf_filter_coeff370_b), 
		.rf_filter_coeff371_a(rf_filter_coeff371_a), 
		.rf_filter_coeff371_b(rf_filter_coeff371_b), 
		.rf_filter_coeff372_a(rf_filter_coeff372_a), 
		.rf_filter_coeff372_b(rf_filter_coeff372_b), 
		.rf_filter_coeff373_a(rf_filter_coeff373_a), 
		.rf_filter_coeff373_b(rf_filter_coeff373_b), 
		.rf_filter_coeff374_a(rf_filter_coeff374_a), 
		.rf_filter_coeff374_b(rf_filter_coeff374_b), 
		.rf_filter_coeff375_a(rf_filter_coeff375_a), 
		.rf_filter_coeff375_b(rf_filter_coeff375_b), 
		.rf_filter_coeff376_a(rf_filter_coeff376_a), 
		.rf_filter_coeff376_b(rf_filter_coeff376_b), 
		.rf_filter_coeff377_a(rf_filter_coeff377_a), 
		.rf_filter_coeff377_b(rf_filter_coeff377_b), 
		.rf_filter_coeff378_a(rf_filter_coeff378_a), 
		.rf_filter_coeff378_b(rf_filter_coeff378_b), 
		.rf_filter_coeff379_a(rf_filter_coeff379_a), 
		.rf_filter_coeff379_b(rf_filter_coeff379_b), 
		.rf_filter_coeff380_a(rf_filter_coeff380_a), 
		.rf_filter_coeff380_b(rf_filter_coeff380_b), 
		.rf_filter_coeff381_a(rf_filter_coeff381_a), 
		.rf_filter_coeff381_b(rf_filter_coeff381_b), 
		.rf_filter_coeff382_a(rf_filter_coeff382_a), 
		.rf_filter_coeff382_b(rf_filter_coeff382_b), 
		.rf_filter_coeff383_a(rf_filter_coeff383_a), 
		.rf_filter_coeff383_b(rf_filter_coeff383_b), 
		.rf_filter_coeff384_a(rf_filter_coeff384_a), 
		.rf_filter_coeff384_b(rf_filter_coeff384_b), 
		.rf_filter_coeff385_a(rf_filter_coeff385_a), 
		.rf_filter_coeff385_b(rf_filter_coeff385_b), 
		.rf_filter_coeff386_a(rf_filter_coeff386_a), 
		.rf_filter_coeff386_b(rf_filter_coeff386_b), 
		.rf_filter_coeff387_a(rf_filter_coeff387_a), 
		.rf_filter_coeff387_b(rf_filter_coeff387_b), 
		.rf_filter_coeff388_a(rf_filter_coeff388_a), 
		.rf_filter_coeff388_b(rf_filter_coeff388_b), 
		.rf_filter_coeff389_a(rf_filter_coeff389_a), 
		.rf_filter_coeff389_b(rf_filter_coeff389_b), 
		.rf_filter_coeff390_a(rf_filter_coeff390_a), 
		.rf_filter_coeff390_b(rf_filter_coeff390_b), 
		.rf_filter_coeff391_a(rf_filter_coeff391_a), 
		.rf_filter_coeff391_b(rf_filter_coeff391_b), 
		.rf_filter_coeff392_a(rf_filter_coeff392_a), 
		.rf_filter_coeff392_b(rf_filter_coeff392_b), 
		.rf_filter_coeff393_a(rf_filter_coeff393_a), 
		.rf_filter_coeff393_b(rf_filter_coeff393_b), 
		.rf_filter_coeff394_a(rf_filter_coeff394_a), 
		.rf_filter_coeff394_b(rf_filter_coeff394_b), 
		.rf_filter_coeff395_a(rf_filter_coeff395_a), 
		.rf_filter_coeff395_b(rf_filter_coeff395_b), 
		.rf_filter_coeff396_a(rf_filter_coeff396_a), 
		.rf_filter_coeff396_b(rf_filter_coeff396_b), 
		.rf_filter_coeff397_a(rf_filter_coeff397_a), 
		.rf_filter_coeff397_b(rf_filter_coeff397_b), 
		.rf_filter_coeff398_a(rf_filter_coeff398_a), 
		.rf_filter_coeff398_b(rf_filter_coeff398_b), 
		.rf_filter_coeff399_a(rf_filter_coeff399_a), 
		.rf_filter_coeff399_b(rf_filter_coeff399_b), 
		.rf_filter_coeff400_a(rf_filter_coeff400_a), 
		.rf_filter_coeff400_b(rf_filter_coeff400_b), 
		.rf_filter_coeff401_a(rf_filter_coeff401_a), 
		.rf_filter_coeff401_b(rf_filter_coeff401_b), 
		.rf_filter_coeff402_a(rf_filter_coeff402_a), 
		.rf_filter_coeff402_b(rf_filter_coeff402_b), 
		.rf_filter_coeff403_a(rf_filter_coeff403_a), 
		.rf_filter_coeff403_b(rf_filter_coeff403_b), 
		.rf_filter_coeff404_a(rf_filter_coeff404_a), 
		.rf_filter_coeff404_b(rf_filter_coeff404_b), 
		.rf_filter_coeff405_a(rf_filter_coeff405_a), 
		.rf_filter_coeff405_b(rf_filter_coeff405_b), 
		.rf_filter_coeff406_a(rf_filter_coeff406_a), 
		.rf_filter_coeff406_b(rf_filter_coeff406_b), 
		.rf_filter_coeff407_a(rf_filter_coeff407_a), 
		.rf_filter_coeff407_b(rf_filter_coeff407_b), 
		.rf_filter_coeff408_a(rf_filter_coeff408_a), 
		.rf_filter_coeff408_b(rf_filter_coeff408_b), 
		.rf_filter_coeff409_a(rf_filter_coeff409_a), 
		.rf_filter_coeff409_b(rf_filter_coeff409_b), 
		.rf_filter_coeff410_a(rf_filter_coeff410_a), 
		.rf_filter_coeff410_b(rf_filter_coeff410_b), 
		.rf_filter_coeff411_a(rf_filter_coeff411_a), 
		.rf_filter_coeff411_b(rf_filter_coeff411_b), 
		.rf_filter_coeff412_a(rf_filter_coeff412_a), 
		.rf_filter_coeff412_b(rf_filter_coeff412_b), 
		.rf_filter_coeff413_a(rf_filter_coeff413_a), 
		.rf_filter_coeff413_b(rf_filter_coeff413_b), 
		.rf_filter_coeff414_a(rf_filter_coeff414_a), 
		.rf_filter_coeff414_b(rf_filter_coeff414_b), 
		.rf_filter_coeff415_a(rf_filter_coeff415_a), 
		.rf_filter_coeff415_b(rf_filter_coeff415_b), 
		.rf_filter_coeff416_a(rf_filter_coeff416_a), 
		.rf_filter_coeff416_b(rf_filter_coeff416_b), 
		.rf_filter_coeff417_a(rf_filter_coeff417_a), 
		.rf_filter_coeff417_b(rf_filter_coeff417_b), 
		.rf_filter_coeff418_a(rf_filter_coeff418_a), 
		.rf_filter_coeff418_b(rf_filter_coeff418_b), 
		.rf_filter_coeff419_a(rf_filter_coeff419_a), 
		.rf_filter_coeff419_b(rf_filter_coeff419_b), 
		.rf_filter_coeff420_a(rf_filter_coeff420_a), 
		.rf_filter_coeff420_b(rf_filter_coeff420_b), 
		.rf_filter_coeff421_a(rf_filter_coeff421_a), 
		.rf_filter_coeff421_b(rf_filter_coeff421_b), 
		.rf_filter_coeff422_a(rf_filter_coeff422_a), 
		.rf_filter_coeff422_b(rf_filter_coeff422_b), 
		.rf_filter_coeff423_a(rf_filter_coeff423_a), 
		.rf_filter_coeff423_b(rf_filter_coeff423_b), 
		.rf_filter_coeff424_a(rf_filter_coeff424_a), 
		.rf_filter_coeff424_b(rf_filter_coeff424_b), 
		.rf_filter_coeff425_a(rf_filter_coeff425_a), 
		.rf_filter_coeff425_b(rf_filter_coeff425_b), 
		.rf_filter_coeff426_a(rf_filter_coeff426_a), 
		.rf_filter_coeff426_b(rf_filter_coeff426_b), 
		.rf_filter_coeff427_a(rf_filter_coeff427_a), 
		.rf_filter_coeff427_b(rf_filter_coeff427_b), 
		.rf_filter_coeff428_a(rf_filter_coeff428_a), 
		.rf_filter_coeff428_b(rf_filter_coeff428_b), 
		.rf_filter_coeff429_a(rf_filter_coeff429_a), 
		.rf_filter_coeff429_b(rf_filter_coeff429_b), 
		.rf_filter_coeff430_a(rf_filter_coeff430_a), 
		.rf_filter_coeff430_b(rf_filter_coeff430_b), 
		.rf_filter_coeff431_a(rf_filter_coeff431_a), 
		.rf_filter_coeff431_b(rf_filter_coeff431_b), 
		.rf_filter_coeff432_a(rf_filter_coeff432_a), 
		.rf_filter_coeff432_b(rf_filter_coeff432_b), 
		.rf_filter_coeff433_a(rf_filter_coeff433_a), 
		.rf_filter_coeff433_b(rf_filter_coeff433_b), 
		.rf_filter_coeff434_a(rf_filter_coeff434_a), 
		.rf_filter_coeff434_b(rf_filter_coeff434_b), 
		.rf_filter_coeff435_a(rf_filter_coeff435_a), 
		.rf_filter_coeff435_b(rf_filter_coeff435_b), 
		.rf_filter_coeff436_a(rf_filter_coeff436_a), 
		.rf_filter_coeff436_b(rf_filter_coeff436_b), 
		.rf_filter_coeff437_a(rf_filter_coeff437_a), 
		.rf_filter_coeff437_b(rf_filter_coeff437_b), 
		.rf_filter_coeff438_a(rf_filter_coeff438_a), 
		.rf_filter_coeff438_b(rf_filter_coeff438_b), 
		.rf_filter_coeff439_a(rf_filter_coeff439_a), 
		.rf_filter_coeff439_b(rf_filter_coeff439_b), 
		.rf_filter_coeff440_a(rf_filter_coeff440_a), 
		.rf_filter_coeff440_b(rf_filter_coeff440_b), 
		.rf_filter_coeff441_a(rf_filter_coeff441_a), 
		.rf_filter_coeff441_b(rf_filter_coeff441_b), 
		.rf_filter_coeff442_a(rf_filter_coeff442_a), 
		.rf_filter_coeff442_b(rf_filter_coeff442_b), 
		.rf_filter_coeff443_a(rf_filter_coeff443_a), 
		.rf_filter_coeff443_b(rf_filter_coeff443_b), 
		.rf_filter_coeff444_a(rf_filter_coeff444_a), 
		.rf_filter_coeff444_b(rf_filter_coeff444_b), 
		.rf_filter_coeff445_a(rf_filter_coeff445_a), 
		.rf_filter_coeff445_b(rf_filter_coeff445_b), 
		.rf_filter_coeff446_a(rf_filter_coeff446_a), 
		.rf_filter_coeff446_b(rf_filter_coeff446_b), 
		.rf_filter_coeff447_a(rf_filter_coeff447_a), 
		.rf_filter_coeff447_b(rf_filter_coeff447_b), 
		.rf_filter_coeff448_a(rf_filter_coeff448_a), 
		.rf_filter_coeff448_b(rf_filter_coeff448_b), 
		.rf_filter_coeff449_a(rf_filter_coeff449_a), 
		.rf_filter_coeff449_b(rf_filter_coeff449_b), 
		.rf_filter_coeff450_a(rf_filter_coeff450_a), 
		.rf_filter_coeff450_b(rf_filter_coeff450_b), 
		.rf_filter_coeff451_a(rf_filter_coeff451_a), 
		.rf_filter_coeff451_b(rf_filter_coeff451_b), 
		.rf_filter_coeff452_a(rf_filter_coeff452_a), 
		.rf_filter_coeff452_b(rf_filter_coeff452_b), 
		.rf_filter_coeff453_a(rf_filter_coeff453_a), 
		.rf_filter_coeff453_b(rf_filter_coeff453_b), 
		.rf_filter_coeff454_a(rf_filter_coeff454_a), 
		.rf_filter_coeff454_b(rf_filter_coeff454_b), 
		.rf_filter_coeff455_a(rf_filter_coeff455_a), 
		.rf_filter_coeff455_b(rf_filter_coeff455_b), 
		.rf_filter_coeff456_a(rf_filter_coeff456_a), 
		.rf_filter_coeff456_b(rf_filter_coeff456_b), 
		.rf_filter_coeff457_a(rf_filter_coeff457_a), 
		.rf_filter_coeff457_b(rf_filter_coeff457_b), 
		.rf_filter_coeff458_a(rf_filter_coeff458_a), 
		.rf_filter_coeff458_b(rf_filter_coeff458_b), 
		.rf_filter_coeff459_a(rf_filter_coeff459_a), 
		.rf_filter_coeff459_b(rf_filter_coeff459_b), 
		.rf_filter_coeff460_a(rf_filter_coeff460_a), 
		.rf_filter_coeff460_b(rf_filter_coeff460_b), 
		.rf_filter_coeff461_a(rf_filter_coeff461_a), 
		.rf_filter_coeff461_b(rf_filter_coeff461_b), 
		.rf_filter_coeff462_a(rf_filter_coeff462_a), 
		.rf_filter_coeff462_b(rf_filter_coeff462_b), 
		.rf_filter_coeff463_a(rf_filter_coeff463_a), 
		.rf_filter_coeff463_b(rf_filter_coeff463_b), 
		.rf_filter_coeff464_a(rf_filter_coeff464_a), 
		.rf_filter_coeff464_b(rf_filter_coeff464_b), 
		.rf_filter_coeff465_a(rf_filter_coeff465_a), 
		.rf_filter_coeff465_b(rf_filter_coeff465_b), 
		.rf_filter_coeff466_a(rf_filter_coeff466_a), 
		.rf_filter_coeff466_b(rf_filter_coeff466_b), 
		.rf_filter_coeff467_a(rf_filter_coeff467_a), 
		.rf_filter_coeff467_b(rf_filter_coeff467_b), 
		.rf_filter_coeff468_a(rf_filter_coeff468_a), 
		.rf_filter_coeff468_b(rf_filter_coeff468_b), 
		.rf_filter_coeff469_a(rf_filter_coeff469_a), 
		.rf_filter_coeff469_b(rf_filter_coeff469_b), 
		.rf_filter_coeff470_a(rf_filter_coeff470_a), 
		.rf_filter_coeff470_b(rf_filter_coeff470_b), 
		.rf_filter_coeff471_a(rf_filter_coeff471_a), 
		.rf_filter_coeff471_b(rf_filter_coeff471_b), 
		.rf_filter_coeff472_a(rf_filter_coeff472_a), 
		.rf_filter_coeff472_b(rf_filter_coeff472_b), 
		.rf_filter_coeff473_a(rf_filter_coeff473_a), 
		.rf_filter_coeff473_b(rf_filter_coeff473_b), 
		.rf_filter_coeff474_a(rf_filter_coeff474_a), 
		.rf_filter_coeff474_b(rf_filter_coeff474_b), 
		.rf_filter_coeff475_a(rf_filter_coeff475_a), 
		.rf_filter_coeff475_b(rf_filter_coeff475_b), 
		.rf_filter_coeff476_a(rf_filter_coeff476_a), 
		.rf_filter_coeff476_b(rf_filter_coeff476_b), 
		.rf_filter_coeff477_a(rf_filter_coeff477_a), 
		.rf_filter_coeff477_b(rf_filter_coeff477_b), 
		.rf_filter_coeff478_a(rf_filter_coeff478_a), 
		.rf_filter_coeff478_b(rf_filter_coeff478_b), 
		.rf_filter_coeff479_a(rf_filter_coeff479_a), 
		.rf_filter_coeff479_b(rf_filter_coeff479_b), 
		.rf_filter_coeff480_a(rf_filter_coeff480_a), 
		.rf_filter_coeff480_b(rf_filter_coeff480_b), 
		.rf_filter_coeff481_a(rf_filter_coeff481_a), 
		.rf_filter_coeff481_b(rf_filter_coeff481_b), 
		.rf_filter_coeff482_a(rf_filter_coeff482_a), 
		.rf_filter_coeff482_b(rf_filter_coeff482_b), 
		.rf_filter_coeff483_a(rf_filter_coeff483_a), 
		.rf_filter_coeff483_b(rf_filter_coeff483_b), 
		.rf_filter_coeff484_a(rf_filter_coeff484_a), 
		.rf_filter_coeff484_b(rf_filter_coeff484_b), 
		.rf_filter_coeff485_a(rf_filter_coeff485_a), 
		.rf_filter_coeff485_b(rf_filter_coeff485_b), 
		.rf_filter_coeff486_a(rf_filter_coeff486_a), 
		.rf_filter_coeff486_b(rf_filter_coeff486_b), 
		.rf_filter_coeff487_a(rf_filter_coeff487_a), 
		.rf_filter_coeff487_b(rf_filter_coeff487_b), 
		.rf_filter_coeff488_a(rf_filter_coeff488_a), 
		.rf_filter_coeff488_b(rf_filter_coeff488_b), 
		.rf_filter_coeff489_a(rf_filter_coeff489_a), 
		.rf_filter_coeff489_b(rf_filter_coeff489_b), 
		.rf_filter_coeff490_a(rf_filter_coeff490_a), 
		.rf_filter_coeff490_b(rf_filter_coeff490_b), 
		.rf_filter_coeff491_a(rf_filter_coeff491_a), 
		.rf_filter_coeff491_b(rf_filter_coeff491_b), 
		.rf_filter_coeff492_a(rf_filter_coeff492_a), 
		.rf_filter_coeff492_b(rf_filter_coeff492_b), 
		.rf_filter_coeff493_a(rf_filter_coeff493_a), 
		.rf_filter_coeff493_b(rf_filter_coeff493_b), 
		.rf_filter_coeff494_a(rf_filter_coeff494_a), 
		.rf_filter_coeff494_b(rf_filter_coeff494_b), 
		.rf_filter_coeff495_a(rf_filter_coeff495_a), 
		.rf_filter_coeff495_b(rf_filter_coeff495_b), 
		.rf_filter_coeff496_a(rf_filter_coeff496_a), 
		.rf_filter_coeff496_b(rf_filter_coeff496_b), 
		.rf_filter_coeff497_a(rf_filter_coeff497_a), 
		.rf_filter_coeff497_b(rf_filter_coeff497_b), 
		.rf_filter_coeff498_a(rf_filter_coeff498_a), 
		.rf_filter_coeff498_b(rf_filter_coeff498_b), 
		.rf_filter_coeff499_a(rf_filter_coeff499_a), 
		.rf_filter_coeff499_b(rf_filter_coeff499_b), 
		.rf_filter_coeff500_a(rf_filter_coeff500_a), 
		.rf_filter_coeff500_b(rf_filter_coeff500_b), 
		.rf_filter_coeff501_a(rf_filter_coeff501_a), 
		.rf_filter_coeff501_b(rf_filter_coeff501_b), 
		.rf_filter_coeff502_a(rf_filter_coeff502_a), 
		.rf_filter_coeff502_b(rf_filter_coeff502_b), 
		.rf_filter_coeff503_a(rf_filter_coeff503_a), 
		.rf_filter_coeff503_b(rf_filter_coeff503_b), 
		.rf_filter_coeff504_a(rf_filter_coeff504_a), 
		.rf_filter_coeff504_b(rf_filter_coeff504_b), 
		.rf_filter_coeff505_a(rf_filter_coeff505_a), 
		.rf_filter_coeff505_b(rf_filter_coeff505_b), 
		.rf_filter_coeff506_a(rf_filter_coeff506_a), 
		.rf_filter_coeff506_b(rf_filter_coeff506_b), 
		.rf_filter_coeff507_a(rf_filter_coeff507_a), 
		.rf_filter_coeff507_b(rf_filter_coeff507_b), 
		.rf_filter_coeff508_a(rf_filter_coeff508_a), 
		.rf_filter_coeff508_b(rf_filter_coeff508_b), 
		.rf_filter_coeff509_a(rf_filter_coeff509_a), 
		.rf_filter_coeff509_b(rf_filter_coeff509_b), 
		.rf_filter_coeff510_a(rf_filter_coeff510_a), 
		.rf_filter_coeff510_b(rf_filter_coeff510_b), 
		.rf_filter_coeff511_a(rf_filter_coeff511_a), 
		.rf_filter_coeff511_b(rf_filter_coeff511_b)
	);

	initial begin
		// Initialize Inputs
		clk = 0;
		rstb = 0;
		//filt_input_data = 32'b00000000000000000100000000000000;
		filt_input_data = 32'h21AB84C2;
		aud_in_rts = 0;
		aud_out_rtr = 0;
		rf_filter_shift = 0;
		rf_filter_clip_en = 0;
		trig_filter_ovf_flag_clear = 0;
		rf_filter_coeff0_a = 1'b1;
		rf_filter_coeff0_b = 0;
		rf_filter_coeff1_a = 0;
		rf_filter_coeff1_b = 0;
		rf_filter_coeff2_a = 0;
		rf_filter_coeff2_b = 0;
		rf_filter_coeff3_a = 0;
		rf_filter_coeff3_b = 0;
		rf_filter_coeff4_a = 0;
		rf_filter_coeff4_b = 0;
		rf_filter_coeff5_a = 0;
		rf_filter_coeff5_b = 0;
		rf_filter_coeff6_a = 0;
		rf_filter_coeff6_b = 0;
		rf_filter_coeff7_a = 0;
		rf_filter_coeff7_b = 0;
		rf_filter_coeff8_a = 0;
		rf_filter_coeff8_b = 0;
		rf_filter_coeff9_a = 0;
		rf_filter_coeff9_b = 0;
		rf_filter_coeff10_a = 0;
		rf_filter_coeff10_b = 0;
		rf_filter_coeff11_a = 0;
		rf_filter_coeff11_b = 0;
		rf_filter_coeff12_a = 0;
		rf_filter_coeff12_b = 0;
		rf_filter_coeff13_a = 0;
		rf_filter_coeff13_b = 0;
		rf_filter_coeff14_a = 0;
		rf_filter_coeff14_b = 0;
		rf_filter_coeff15_a = 0;
		rf_filter_coeff15_b = 0;
		rf_filter_coeff16_a = 0;
		rf_filter_coeff16_b = 0;
		rf_filter_coeff17_a = 0;
		rf_filter_coeff17_b = 0;
		rf_filter_coeff18_a = 0;
		rf_filter_coeff18_b = 0;
		rf_filter_coeff19_a = 0;
		rf_filter_coeff19_b = 0;
		rf_filter_coeff20_a = 0;
		rf_filter_coeff20_b = 0;
		rf_filter_coeff21_a = 0;
		rf_filter_coeff21_b = 0;
		rf_filter_coeff22_a = 0;
		rf_filter_coeff22_b = 0;
		rf_filter_coeff23_a = 0;
		rf_filter_coeff23_b = 0;
		rf_filter_coeff24_a = 0;
		rf_filter_coeff24_b = 0;
		rf_filter_coeff25_a = 0;
		rf_filter_coeff25_b = 0;
		rf_filter_coeff26_a = 0;
		rf_filter_coeff26_b = 0;
		rf_filter_coeff27_a = 0;
		rf_filter_coeff27_b = 0;
		rf_filter_coeff28_a = 0;
		rf_filter_coeff28_b = 0;
		rf_filter_coeff29_a = 0;
		rf_filter_coeff29_b = 0;
		rf_filter_coeff30_a = 0;
		rf_filter_coeff30_b = 0;
		rf_filter_coeff31_a = 0;
		rf_filter_coeff31_b = 0;
		rf_filter_coeff32_a = 0;
		rf_filter_coeff32_b = 0;
		rf_filter_coeff33_a = 0;
		rf_filter_coeff33_b = 0;
		rf_filter_coeff34_a = 0;
		rf_filter_coeff34_b = 0;
		rf_filter_coeff35_a = 0;
		rf_filter_coeff35_b = 0;
		rf_filter_coeff36_a = 0;
		rf_filter_coeff36_b = 0;
		rf_filter_coeff37_a = 0;
		rf_filter_coeff37_b = 0;
		rf_filter_coeff38_a = 0;
		rf_filter_coeff38_b = 0;
		rf_filter_coeff39_a = 0;
		rf_filter_coeff39_b = 0;
		rf_filter_coeff40_a = 0;
		rf_filter_coeff40_b = 0;
		rf_filter_coeff41_a = 0;
		rf_filter_coeff41_b = 0;
		rf_filter_coeff42_a = 0;
		rf_filter_coeff42_b = 0;
		rf_filter_coeff43_a = 0;
		rf_filter_coeff43_b = 0;
		rf_filter_coeff44_a = 0;
		rf_filter_coeff44_b = 0;
		rf_filter_coeff45_a = 0;
		rf_filter_coeff45_b = 0;
		rf_filter_coeff46_a = 0;
		rf_filter_coeff46_b = 0;
		rf_filter_coeff47_a = 0;
		rf_filter_coeff47_b = 0;
		rf_filter_coeff48_a = 0;
		rf_filter_coeff48_b = 0;
		rf_filter_coeff49_a = 0;
		rf_filter_coeff49_b = 0;
		rf_filter_coeff50_a = 0;
		rf_filter_coeff50_b = 0;
		rf_filter_coeff51_a = 0;
		rf_filter_coeff51_b = 0;
		rf_filter_coeff52_a = 0;
		rf_filter_coeff52_b = 0;
		rf_filter_coeff53_a = 0;
		rf_filter_coeff53_b = 0;
		rf_filter_coeff54_a = 0;
		rf_filter_coeff54_b = 0;
		rf_filter_coeff55_a = 0;
		rf_filter_coeff55_b = 0;
		rf_filter_coeff56_a = 0;
		rf_filter_coeff56_b = 0;
		rf_filter_coeff57_a = 0;
		rf_filter_coeff57_b = 0;
		rf_filter_coeff58_a = 0;
		rf_filter_coeff58_b = 0;
		rf_filter_coeff59_a = 0;
		rf_filter_coeff59_b = 0;
		rf_filter_coeff60_a = 0;
		rf_filter_coeff60_b = 0;
		rf_filter_coeff61_a = 0;
		rf_filter_coeff61_b = 0;
		rf_filter_coeff62_a = 0;
		rf_filter_coeff62_b = 0;
		rf_filter_coeff63_a = 0;
		rf_filter_coeff63_b = 0;
		rf_filter_coeff64_a = 0;
		rf_filter_coeff64_b = 0;
		rf_filter_coeff65_a = 0;
		rf_filter_coeff65_b = 0;
		rf_filter_coeff66_a = 0;
		rf_filter_coeff66_b = 0;
		rf_filter_coeff67_a = 0;
		rf_filter_coeff67_b = 0;
		rf_filter_coeff68_a = 0;
		rf_filter_coeff68_b = 0;
		rf_filter_coeff69_a = 0;
		rf_filter_coeff69_b = 0;
		rf_filter_coeff70_a = 0;
		rf_filter_coeff70_b = 0;
		rf_filter_coeff71_a = 0;
		rf_filter_coeff71_b = 0;
		rf_filter_coeff72_a = 0;
		rf_filter_coeff72_b = 0;
		rf_filter_coeff73_a = 0;
		rf_filter_coeff73_b = 0;
		rf_filter_coeff74_a = 0;
		rf_filter_coeff74_b = 0;
		rf_filter_coeff75_a = 0;
		rf_filter_coeff75_b = 0;
		rf_filter_coeff76_a = 0;
		rf_filter_coeff76_b = 0;
		rf_filter_coeff77_a = 0;
		rf_filter_coeff77_b = 0;
		rf_filter_coeff78_a = 0;
		rf_filter_coeff78_b = 0;
		rf_filter_coeff79_a = 0;
		rf_filter_coeff79_b = 0;
		rf_filter_coeff80_a = 0;
		rf_filter_coeff80_b = 0;
		rf_filter_coeff81_a = 0;
		rf_filter_coeff81_b = 0;
		rf_filter_coeff82_a = 0;
		rf_filter_coeff82_b = 0;
		rf_filter_coeff83_a = 0;
		rf_filter_coeff83_b = 0;
		rf_filter_coeff84_a = 0;
		rf_filter_coeff84_b = 0;
		rf_filter_coeff85_a = 0;
		rf_filter_coeff85_b = 0;
		rf_filter_coeff86_a = 0;
		rf_filter_coeff86_b = 0;
		rf_filter_coeff87_a = 0;
		rf_filter_coeff87_b = 0;
		rf_filter_coeff88_a = 0;
		rf_filter_coeff88_b = 0;
		rf_filter_coeff89_a = 0;
		rf_filter_coeff89_b = 0;
		rf_filter_coeff90_a = 0;
		rf_filter_coeff90_b = 0;
		rf_filter_coeff91_a = 0;
		rf_filter_coeff91_b = 0;
		rf_filter_coeff92_a = 0;
		rf_filter_coeff92_b = 0;
		rf_filter_coeff93_a = 0;
		rf_filter_coeff93_b = 0;
		rf_filter_coeff94_a = 0;
		rf_filter_coeff94_b = 0;
		rf_filter_coeff95_a = 0;
		rf_filter_coeff95_b = 0;
		rf_filter_coeff96_a = 0;
		rf_filter_coeff96_b = 0;
		rf_filter_coeff97_a = 0;
		rf_filter_coeff97_b = 0;
		rf_filter_coeff98_a = 0;
		rf_filter_coeff98_b = 0;
		rf_filter_coeff99_a = 0;
		rf_filter_coeff99_b = 0;
		rf_filter_coeff100_a = 0;
		rf_filter_coeff100_b = 0;
		rf_filter_coeff101_a = 0;
		rf_filter_coeff101_b = 0;
		rf_filter_coeff102_a = 0;
		rf_filter_coeff102_b = 0;
		rf_filter_coeff103_a = 0;
		rf_filter_coeff103_b = 0;
		rf_filter_coeff104_a = 0;
		rf_filter_coeff104_b = 0;
		rf_filter_coeff105_a = 0;
		rf_filter_coeff105_b = 0;
		rf_filter_coeff106_a = 0;
		rf_filter_coeff106_b = 0;
		rf_filter_coeff107_a = 0;
		rf_filter_coeff107_b = 0;
		rf_filter_coeff108_a = 0;
		rf_filter_coeff108_b = 0;
		rf_filter_coeff109_a = 0;
		rf_filter_coeff109_b = 0;
		rf_filter_coeff110_a = 0;
		rf_filter_coeff110_b = 0;
		rf_filter_coeff111_a = 0;
		rf_filter_coeff111_b = 0;
		rf_filter_coeff112_a = 0;
		rf_filter_coeff112_b = 0;
		rf_filter_coeff113_a = 0;
		rf_filter_coeff113_b = 0;
		rf_filter_coeff114_a = 0;
		rf_filter_coeff114_b = 0;
		rf_filter_coeff115_a = 0;
		rf_filter_coeff115_b = 0;
		rf_filter_coeff116_a = 0;
		rf_filter_coeff116_b = 0;
		rf_filter_coeff117_a = 0;
		rf_filter_coeff117_b = 0;
		rf_filter_coeff118_a = 0;
		rf_filter_coeff118_b = 0;
		rf_filter_coeff119_a = 0;
		rf_filter_coeff119_b = 0;
		rf_filter_coeff120_a = 0;
		rf_filter_coeff120_b = 0;
		rf_filter_coeff121_a = 0;
		rf_filter_coeff121_b = 0;
		rf_filter_coeff122_a = 0;
		rf_filter_coeff122_b = 0;
		rf_filter_coeff123_a = 0;
		rf_filter_coeff123_b = 0;
		rf_filter_coeff124_a = 0;
		rf_filter_coeff124_b = 0;
		rf_filter_coeff125_a = 0;
		rf_filter_coeff125_b = 0;
		rf_filter_coeff126_a = 0;
		rf_filter_coeff126_b = 0;
		rf_filter_coeff127_a = 0;
		rf_filter_coeff127_b = 0;
		rf_filter_coeff128_a = 0;
		rf_filter_coeff128_b = 0;
		rf_filter_coeff129_a = 0;
		rf_filter_coeff129_b = 0;
		rf_filter_coeff130_a = 0;
		rf_filter_coeff130_b = 0;
		rf_filter_coeff131_a = 0;
		rf_filter_coeff131_b = 0;
		rf_filter_coeff132_a = 0;
		rf_filter_coeff132_b = 0;
		rf_filter_coeff133_a = 0;
		rf_filter_coeff133_b = 0;
		rf_filter_coeff134_a = 0;
		rf_filter_coeff134_b = 0;
		rf_filter_coeff135_a = 0;
		rf_filter_coeff135_b = 0;
		rf_filter_coeff136_a = 0;
		rf_filter_coeff136_b = 0;
		rf_filter_coeff137_a = 0;
		rf_filter_coeff137_b = 0;
		rf_filter_coeff138_a = 0;
		rf_filter_coeff138_b = 0;
		rf_filter_coeff139_a = 0;
		rf_filter_coeff139_b = 0;
		rf_filter_coeff140_a = 0;
		rf_filter_coeff140_b = 0;
		rf_filter_coeff141_a = 0;
		rf_filter_coeff141_b = 0;
		rf_filter_coeff142_a = 0;
		rf_filter_coeff142_b = 0;
		rf_filter_coeff143_a = 0;
		rf_filter_coeff143_b = 0;
		rf_filter_coeff144_a = 0;
		rf_filter_coeff144_b = 0;
		rf_filter_coeff145_a = 0;
		rf_filter_coeff145_b = 0;
		rf_filter_coeff146_a = 0;
		rf_filter_coeff146_b = 0;
		rf_filter_coeff147_a = 0;
		rf_filter_coeff147_b = 0;
		rf_filter_coeff148_a = 0;
		rf_filter_coeff148_b = 0;
		rf_filter_coeff149_a = 0;
		rf_filter_coeff149_b = 0;
		rf_filter_coeff150_a = 0;
		rf_filter_coeff150_b = 0;
		rf_filter_coeff151_a = 0;
		rf_filter_coeff151_b = 0;
		rf_filter_coeff152_a = 0;
		rf_filter_coeff152_b = 0;
		rf_filter_coeff153_a = 0;
		rf_filter_coeff153_b = 0;
		rf_filter_coeff154_a = 0;
		rf_filter_coeff154_b = 0;
		rf_filter_coeff155_a = 0;
		rf_filter_coeff155_b = 0;
		rf_filter_coeff156_a = 0;
		rf_filter_coeff156_b = 0;
		rf_filter_coeff157_a = 0;
		rf_filter_coeff157_b = 0;
		rf_filter_coeff158_a = 0;
		rf_filter_coeff158_b = 0;
		rf_filter_coeff159_a = 0;
		rf_filter_coeff159_b = 0;
		rf_filter_coeff160_a = 0;
		rf_filter_coeff160_b = 0;
		rf_filter_coeff161_a = 0;
		rf_filter_coeff161_b = 0;
		rf_filter_coeff162_a = 0;
		rf_filter_coeff162_b = 0;
		rf_filter_coeff163_a = 0;
		rf_filter_coeff163_b = 0;
		rf_filter_coeff164_a = 0;
		rf_filter_coeff164_b = 0;
		rf_filter_coeff165_a = 0;
		rf_filter_coeff165_b = 0;
		rf_filter_coeff166_a = 0;
		rf_filter_coeff166_b = 0;
		rf_filter_coeff167_a = 0;
		rf_filter_coeff167_b = 0;
		rf_filter_coeff168_a = 0;
		rf_filter_coeff168_b = 0;
		rf_filter_coeff169_a = 0;
		rf_filter_coeff169_b = 0;
		rf_filter_coeff170_a = 0;
		rf_filter_coeff170_b = 0;
		rf_filter_coeff171_a = 0;
		rf_filter_coeff171_b = 0;
		rf_filter_coeff172_a = 0;
		rf_filter_coeff172_b = 0;
		rf_filter_coeff173_a = 0;
		rf_filter_coeff173_b = 0;
		rf_filter_coeff174_a = 0;
		rf_filter_coeff174_b = 0;
		rf_filter_coeff175_a = 0;
		rf_filter_coeff175_b = 0;
		rf_filter_coeff176_a = 0;
		rf_filter_coeff176_b = 0;
		rf_filter_coeff177_a = 0;
		rf_filter_coeff177_b = 0;
		rf_filter_coeff178_a = 0;
		rf_filter_coeff178_b = 0;
		rf_filter_coeff179_a = 0;
		rf_filter_coeff179_b = 0;
		rf_filter_coeff180_a = 0;
		rf_filter_coeff180_b = 0;
		rf_filter_coeff181_a = 0;
		rf_filter_coeff181_b = 0;
		rf_filter_coeff182_a = 0;
		rf_filter_coeff182_b = 0;
		rf_filter_coeff183_a = 0;
		rf_filter_coeff183_b = 0;
		rf_filter_coeff184_a = 0;
		rf_filter_coeff184_b = 0;
		rf_filter_coeff185_a = 0;
		rf_filter_coeff185_b = 0;
		rf_filter_coeff186_a = 0;
		rf_filter_coeff186_b = 0;
		rf_filter_coeff187_a = 0;
		rf_filter_coeff187_b = 0;
		rf_filter_coeff188_a = 0;
		rf_filter_coeff188_b = 0;
		rf_filter_coeff189_a = 0;
		rf_filter_coeff189_b = 0;
		rf_filter_coeff190_a = 0;
		rf_filter_coeff190_b = 0;
		rf_filter_coeff191_a = 0;
		rf_filter_coeff191_b = 0;
		rf_filter_coeff192_a = 0;
		rf_filter_coeff192_b = 0;
		rf_filter_coeff193_a = 0;
		rf_filter_coeff193_b = 0;
		rf_filter_coeff194_a = 0;
		rf_filter_coeff194_b = 0;
		rf_filter_coeff195_a = 0;
		rf_filter_coeff195_b = 0;
		rf_filter_coeff196_a = 0;
		rf_filter_coeff196_b = 0;
		rf_filter_coeff197_a = 0;
		rf_filter_coeff197_b = 0;
		rf_filter_coeff198_a = 0;
		rf_filter_coeff198_b = 0;
		rf_filter_coeff199_a = 0;
		rf_filter_coeff199_b = 0;
		rf_filter_coeff200_a = 0;
		rf_filter_coeff200_b = 0;
		rf_filter_coeff201_a = 0;
		rf_filter_coeff201_b = 0;
		rf_filter_coeff202_a = 0;
		rf_filter_coeff202_b = 0;
		rf_filter_coeff203_a = 0;
		rf_filter_coeff203_b = 0;
		rf_filter_coeff204_a = 0;
		rf_filter_coeff204_b = 0;
		rf_filter_coeff205_a = 0;
		rf_filter_coeff205_b = 0;
		rf_filter_coeff206_a = 0;
		rf_filter_coeff206_b = 0;
		rf_filter_coeff207_a = 0;
		rf_filter_coeff207_b = 0;
		rf_filter_coeff208_a = 0;
		rf_filter_coeff208_b = 0;
		rf_filter_coeff209_a = 0;
		rf_filter_coeff209_b = 0;
		rf_filter_coeff210_a = 0;
		rf_filter_coeff210_b = 0;
		rf_filter_coeff211_a = 0;
		rf_filter_coeff211_b = 0;
		rf_filter_coeff212_a = 0;
		rf_filter_coeff212_b = 0;
		rf_filter_coeff213_a = 0;
		rf_filter_coeff213_b = 0;
		rf_filter_coeff214_a = 0;
		rf_filter_coeff214_b = 0;
		rf_filter_coeff215_a = 0;
		rf_filter_coeff215_b = 0;
		rf_filter_coeff216_a = 0;
		rf_filter_coeff216_b = 0;
		rf_filter_coeff217_a = 0;
		rf_filter_coeff217_b = 0;
		rf_filter_coeff218_a = 0;
		rf_filter_coeff218_b = 0;
		rf_filter_coeff219_a = 0;
		rf_filter_coeff219_b = 0;
		rf_filter_coeff220_a = 0;
		rf_filter_coeff220_b = 0;
		rf_filter_coeff221_a = 0;
		rf_filter_coeff221_b = 0;
		rf_filter_coeff222_a = 0;
		rf_filter_coeff222_b = 0;
		rf_filter_coeff223_a = 0;
		rf_filter_coeff223_b = 0;
		rf_filter_coeff224_a = 0;
		rf_filter_coeff224_b = 0;
		rf_filter_coeff225_a = 0;
		rf_filter_coeff225_b = 0;
		rf_filter_coeff226_a = 0;
		rf_filter_coeff226_b = 0;
		rf_filter_coeff227_a = 0;
		rf_filter_coeff227_b = 0;
		rf_filter_coeff228_a = 0;
		rf_filter_coeff228_b = 0;
		rf_filter_coeff229_a = 0;
		rf_filter_coeff229_b = 0;
		rf_filter_coeff230_a = 0;
		rf_filter_coeff230_b = 0;
		rf_filter_coeff231_a = 0;
		rf_filter_coeff231_b = 0;
		rf_filter_coeff232_a = 0;
		rf_filter_coeff232_b = 0;
		rf_filter_coeff233_a = 0;
		rf_filter_coeff233_b = 0;
		rf_filter_coeff234_a = 0;
		rf_filter_coeff234_b = 0;
		rf_filter_coeff235_a = 0;
		rf_filter_coeff235_b = 0;
		rf_filter_coeff236_a = 0;
		rf_filter_coeff236_b = 0;
		rf_filter_coeff237_a = 0;
		rf_filter_coeff237_b = 0;
		rf_filter_coeff238_a = 0;
		rf_filter_coeff238_b = 0;
		rf_filter_coeff239_a = 0;
		rf_filter_coeff239_b = 0;
		rf_filter_coeff240_a = 0;
		rf_filter_coeff240_b = 0;
		rf_filter_coeff241_a = 0;
		rf_filter_coeff241_b = 0;
		rf_filter_coeff242_a = 0;
		rf_filter_coeff242_b = 0;
		rf_filter_coeff243_a = 0;
		rf_filter_coeff243_b = 0;
		rf_filter_coeff244_a = 0;
		rf_filter_coeff244_b = 0;
		rf_filter_coeff245_a = 0;
		rf_filter_coeff245_b = 0;
		rf_filter_coeff246_a = 0;
		rf_filter_coeff246_b = 0;
		rf_filter_coeff247_a = 0;
		rf_filter_coeff247_b = 0;
		rf_filter_coeff248_a = 0;
		rf_filter_coeff248_b = 0;
		rf_filter_coeff249_a = 0;
		rf_filter_coeff249_b = 0;
		rf_filter_coeff250_a = 0;
		rf_filter_coeff250_b = 0;
		rf_filter_coeff251_a = 0;
		rf_filter_coeff251_b = 0;
		rf_filter_coeff252_a = 0;
		rf_filter_coeff252_b = 0;
		rf_filter_coeff253_a = 0;
		rf_filter_coeff253_b = 0;
		rf_filter_coeff254_a = 0;
		rf_filter_coeff254_b = 0;
		rf_filter_coeff255_a = 0;
		rf_filter_coeff255_b = 0;
		rf_filter_coeff256_a = 0;
		rf_filter_coeff256_b = 0;
		rf_filter_coeff257_a = 0;
		rf_filter_coeff257_b = 0;
		rf_filter_coeff258_a = 0;
		rf_filter_coeff258_b = 0;
		rf_filter_coeff259_a = 0;
		rf_filter_coeff259_b = 0;
		rf_filter_coeff260_a = 0;
		rf_filter_coeff260_b = 0;
		rf_filter_coeff261_a = 0;
		rf_filter_coeff261_b = 0;
		rf_filter_coeff262_a = 0;
		rf_filter_coeff262_b = 0;
		rf_filter_coeff263_a = 0;
		rf_filter_coeff263_b = 0;
		rf_filter_coeff264_a = 0;
		rf_filter_coeff264_b = 0;
		rf_filter_coeff265_a = 0;
		rf_filter_coeff265_b = 0;
		rf_filter_coeff266_a = 0;
		rf_filter_coeff266_b = 0;
		rf_filter_coeff267_a = 0;
		rf_filter_coeff267_b = 0;
		rf_filter_coeff268_a = 0;
		rf_filter_coeff268_b = 0;
		rf_filter_coeff269_a = 0;
		rf_filter_coeff269_b = 0;
		rf_filter_coeff270_a = 0;
		rf_filter_coeff270_b = 0;
		rf_filter_coeff271_a = 0;
		rf_filter_coeff271_b = 0;
		rf_filter_coeff272_a = 0;
		rf_filter_coeff272_b = 0;
		rf_filter_coeff273_a = 0;
		rf_filter_coeff273_b = 0;
		rf_filter_coeff274_a = 0;
		rf_filter_coeff274_b = 0;
		rf_filter_coeff275_a = 0;
		rf_filter_coeff275_b = 0;
		rf_filter_coeff276_a = 0;
		rf_filter_coeff276_b = 0;
		rf_filter_coeff277_a = 0;
		rf_filter_coeff277_b = 0;
		rf_filter_coeff278_a = 0;
		rf_filter_coeff278_b = 0;
		rf_filter_coeff279_a = 0;
		rf_filter_coeff279_b = 0;
		rf_filter_coeff280_a = 0;
		rf_filter_coeff280_b = 0;
		rf_filter_coeff281_a = 0;
		rf_filter_coeff281_b = 0;
		rf_filter_coeff282_a = 0;
		rf_filter_coeff282_b = 0;
		rf_filter_coeff283_a = 0;
		rf_filter_coeff283_b = 0;
		rf_filter_coeff284_a = 0;
		rf_filter_coeff284_b = 0;
		rf_filter_coeff285_a = 0;
		rf_filter_coeff285_b = 0;
		rf_filter_coeff286_a = 0;
		rf_filter_coeff286_b = 0;
		rf_filter_coeff287_a = 0;
		rf_filter_coeff287_b = 0;
		rf_filter_coeff288_a = 0;
		rf_filter_coeff288_b = 0;
		rf_filter_coeff289_a = 0;
		rf_filter_coeff289_b = 0;
		rf_filter_coeff290_a = 0;
		rf_filter_coeff290_b = 0;
		rf_filter_coeff291_a = 0;
		rf_filter_coeff291_b = 0;
		rf_filter_coeff292_a = 0;
		rf_filter_coeff292_b = 0;
		rf_filter_coeff293_a = 0;
		rf_filter_coeff293_b = 0;
		rf_filter_coeff294_a = 0;
		rf_filter_coeff294_b = 0;
		rf_filter_coeff295_a = 0;
		rf_filter_coeff295_b = 0;
		rf_filter_coeff296_a = 0;
		rf_filter_coeff296_b = 0;
		rf_filter_coeff297_a = 0;
		rf_filter_coeff297_b = 0;
		rf_filter_coeff298_a = 0;
		rf_filter_coeff298_b = 0;
		rf_filter_coeff299_a = 0;
		rf_filter_coeff299_b = 0;
		rf_filter_coeff300_a = 0;
		rf_filter_coeff300_b = 0;
		rf_filter_coeff301_a = 0;
		rf_filter_coeff301_b = 0;
		rf_filter_coeff302_a = 0;
		rf_filter_coeff302_b = 0;
		rf_filter_coeff303_a = 0;
		rf_filter_coeff303_b = 0;
		rf_filter_coeff304_a = 0;
		rf_filter_coeff304_b = 0;
		rf_filter_coeff305_a = 0;
		rf_filter_coeff305_b = 0;
		rf_filter_coeff306_a = 0;
		rf_filter_coeff306_b = 0;
		rf_filter_coeff307_a = 0;
		rf_filter_coeff307_b = 0;
		rf_filter_coeff308_a = 0;
		rf_filter_coeff308_b = 0;
		rf_filter_coeff309_a = 0;
		rf_filter_coeff309_b = 0;
		rf_filter_coeff310_a = 0;
		rf_filter_coeff310_b = 0;
		rf_filter_coeff311_a = 0;
		rf_filter_coeff311_b = 0;
		rf_filter_coeff312_a = 0;
		rf_filter_coeff312_b = 0;
		rf_filter_coeff313_a = 0;
		rf_filter_coeff313_b = 0;
		rf_filter_coeff314_a = 0;
		rf_filter_coeff314_b = 0;
		rf_filter_coeff315_a = 0;
		rf_filter_coeff315_b = 0;
		rf_filter_coeff316_a = 0;
		rf_filter_coeff316_b = 0;
		rf_filter_coeff317_a = 0;
		rf_filter_coeff317_b = 0;
		rf_filter_coeff318_a = 0;
		rf_filter_coeff318_b = 0;
		rf_filter_coeff319_a = 0;
		rf_filter_coeff319_b = 0;
		rf_filter_coeff320_a = 0;
		rf_filter_coeff320_b = 0;
		rf_filter_coeff321_a = 0;
		rf_filter_coeff321_b = 0;
		rf_filter_coeff322_a = 0;
		rf_filter_coeff322_b = 0;
		rf_filter_coeff323_a = 0;
		rf_filter_coeff323_b = 0;
		rf_filter_coeff324_a = 0;
		rf_filter_coeff324_b = 0;
		rf_filter_coeff325_a = 0;
		rf_filter_coeff325_b = 0;
		rf_filter_coeff326_a = 0;
		rf_filter_coeff326_b = 0;
		rf_filter_coeff327_a = 0;
		rf_filter_coeff327_b = 0;
		rf_filter_coeff328_a = 0;
		rf_filter_coeff328_b = 0;
		rf_filter_coeff329_a = 0;
		rf_filter_coeff329_b = 0;
		rf_filter_coeff330_a = 0;
		rf_filter_coeff330_b = 0;
		rf_filter_coeff331_a = 0;
		rf_filter_coeff331_b = 0;
		rf_filter_coeff332_a = 0;
		rf_filter_coeff332_b = 0;
		rf_filter_coeff333_a = 0;
		rf_filter_coeff333_b = 0;
		rf_filter_coeff334_a = 0;
		rf_filter_coeff334_b = 0;
		rf_filter_coeff335_a = 0;
		rf_filter_coeff335_b = 0;
		rf_filter_coeff336_a = 0;
		rf_filter_coeff336_b = 0;
		rf_filter_coeff337_a = 0;
		rf_filter_coeff337_b = 0;
		rf_filter_coeff338_a = 0;
		rf_filter_coeff338_b = 0;
		rf_filter_coeff339_a = 0;
		rf_filter_coeff339_b = 0;
		rf_filter_coeff340_a = 0;
		rf_filter_coeff340_b = 0;
		rf_filter_coeff341_a = 0;
		rf_filter_coeff341_b = 0;
		rf_filter_coeff342_a = 0;
		rf_filter_coeff342_b = 0;
		rf_filter_coeff343_a = 0;
		rf_filter_coeff343_b = 0;
		rf_filter_coeff344_a = 0;
		rf_filter_coeff344_b = 0;
		rf_filter_coeff345_a = 0;
		rf_filter_coeff345_b = 0;
		rf_filter_coeff346_a = 0;
		rf_filter_coeff346_b = 0;
		rf_filter_coeff347_a = 0;
		rf_filter_coeff347_b = 0;
		rf_filter_coeff348_a = 0;
		rf_filter_coeff348_b = 0;
		rf_filter_coeff349_a = 0;
		rf_filter_coeff349_b = 0;
		rf_filter_coeff350_a = 0;
		rf_filter_coeff350_b = 0;
		rf_filter_coeff351_a = 0;
		rf_filter_coeff351_b = 0;
		rf_filter_coeff352_a = 0;
		rf_filter_coeff352_b = 0;
		rf_filter_coeff353_a = 0;
		rf_filter_coeff353_b = 0;
		rf_filter_coeff354_a = 0;
		rf_filter_coeff354_b = 0;
		rf_filter_coeff355_a = 0;
		rf_filter_coeff355_b = 0;
		rf_filter_coeff356_a = 0;
		rf_filter_coeff356_b = 0;
		rf_filter_coeff357_a = 0;
		rf_filter_coeff357_b = 0;
		rf_filter_coeff358_a = 0;
		rf_filter_coeff358_b = 0;
		rf_filter_coeff359_a = 0;
		rf_filter_coeff359_b = 0;
		rf_filter_coeff360_a = 0;
		rf_filter_coeff360_b = 0;
		rf_filter_coeff361_a = 0;
		rf_filter_coeff361_b = 0;
		rf_filter_coeff362_a = 0;
		rf_filter_coeff362_b = 0;
		rf_filter_coeff363_a = 0;
		rf_filter_coeff363_b = 0;
		rf_filter_coeff364_a = 0;
		rf_filter_coeff364_b = 0;
		rf_filter_coeff365_a = 0;
		rf_filter_coeff365_b = 0;
		rf_filter_coeff366_a = 0;
		rf_filter_coeff366_b = 0;
		rf_filter_coeff367_a = 0;
		rf_filter_coeff367_b = 0;
		rf_filter_coeff368_a = 0;
		rf_filter_coeff368_b = 0;
		rf_filter_coeff369_a = 0;
		rf_filter_coeff369_b = 0;
		rf_filter_coeff370_a = 0;
		rf_filter_coeff370_b = 0;
		rf_filter_coeff371_a = 0;
		rf_filter_coeff371_b = 0;
		rf_filter_coeff372_a = 0;
		rf_filter_coeff372_b = 0;
		rf_filter_coeff373_a = 0;
		rf_filter_coeff373_b = 0;
		rf_filter_coeff374_a = 0;
		rf_filter_coeff374_b = 0;
		rf_filter_coeff375_a = 0;
		rf_filter_coeff375_b = 0;
		rf_filter_coeff376_a = 0;
		rf_filter_coeff376_b = 0;
		rf_filter_coeff377_a = 0;
		rf_filter_coeff377_b = 0;
		rf_filter_coeff378_a = 0;
		rf_filter_coeff378_b = 0;
		rf_filter_coeff379_a = 0;
		rf_filter_coeff379_b = 0;
		rf_filter_coeff380_a = 0;
		rf_filter_coeff380_b = 0;
		rf_filter_coeff381_a = 0;
		rf_filter_coeff381_b = 0;
		rf_filter_coeff382_a = 0;
		rf_filter_coeff382_b = 0;
		rf_filter_coeff383_a = 0;
		rf_filter_coeff383_b = 0;
		rf_filter_coeff384_a = 0;
		rf_filter_coeff384_b = 0;
		rf_filter_coeff385_a = 0;
		rf_filter_coeff385_b = 0;
		rf_filter_coeff386_a = 0;
		rf_filter_coeff386_b = 0;
		rf_filter_coeff387_a = 0;
		rf_filter_coeff387_b = 0;
		rf_filter_coeff388_a = 0;
		rf_filter_coeff388_b = 0;
		rf_filter_coeff389_a = 0;
		rf_filter_coeff389_b = 0;
		rf_filter_coeff390_a = 0;
		rf_filter_coeff390_b = 0;
		rf_filter_coeff391_a = 0;
		rf_filter_coeff391_b = 0;
		rf_filter_coeff392_a = 0;
		rf_filter_coeff392_b = 0;
		rf_filter_coeff393_a = 0;
		rf_filter_coeff393_b = 0;
		rf_filter_coeff394_a = 0;
		rf_filter_coeff394_b = 0;
		rf_filter_coeff395_a = 0;
		rf_filter_coeff395_b = 0;
		rf_filter_coeff396_a = 0;
		rf_filter_coeff396_b = 0;
		rf_filter_coeff397_a = 0;
		rf_filter_coeff397_b = 0;
		rf_filter_coeff398_a = 0;
		rf_filter_coeff398_b = 0;
		rf_filter_coeff399_a = 0;
		rf_filter_coeff399_b = 0;
		rf_filter_coeff400_a = 0;
		rf_filter_coeff400_b = 0;
		rf_filter_coeff401_a = 0;
		rf_filter_coeff401_b = 0;
		rf_filter_coeff402_a = 0;
		rf_filter_coeff402_b = 0;
		rf_filter_coeff403_a = 0;
		rf_filter_coeff403_b = 0;
		rf_filter_coeff404_a = 0;
		rf_filter_coeff404_b = 0;
		rf_filter_coeff405_a = 0;
		rf_filter_coeff405_b = 0;
		rf_filter_coeff406_a = 0;
		rf_filter_coeff406_b = 0;
		rf_filter_coeff407_a = 0;
		rf_filter_coeff407_b = 0;
		rf_filter_coeff408_a = 0;
		rf_filter_coeff408_b = 0;
		rf_filter_coeff409_a = 0;
		rf_filter_coeff409_b = 0;
		rf_filter_coeff410_a = 0;
		rf_filter_coeff410_b = 0;
		rf_filter_coeff411_a = 0;
		rf_filter_coeff411_b = 0;
		rf_filter_coeff412_a = 0;
		rf_filter_coeff412_b = 0;
		rf_filter_coeff413_a = 0;
		rf_filter_coeff413_b = 0;
		rf_filter_coeff414_a = 0;
		rf_filter_coeff414_b = 0;
		rf_filter_coeff415_a = 0;
		rf_filter_coeff415_b = 0;
		rf_filter_coeff416_a = 0;
		rf_filter_coeff416_b = 0;
		rf_filter_coeff417_a = 0;
		rf_filter_coeff417_b = 0;
		rf_filter_coeff418_a = 0;
		rf_filter_coeff418_b = 0;
		rf_filter_coeff419_a = 0;
		rf_filter_coeff419_b = 0;
		rf_filter_coeff420_a = 0;
		rf_filter_coeff420_b = 0;
		rf_filter_coeff421_a = 0;
		rf_filter_coeff421_b = 0;
		rf_filter_coeff422_a = 0;
		rf_filter_coeff422_b = 0;
		rf_filter_coeff423_a = 0;
		rf_filter_coeff423_b = 0;
		rf_filter_coeff424_a = 0;
		rf_filter_coeff424_b = 0;
		rf_filter_coeff425_a = 0;
		rf_filter_coeff425_b = 0;
		rf_filter_coeff426_a = 0;
		rf_filter_coeff426_b = 0;
		rf_filter_coeff427_a = 0;
		rf_filter_coeff427_b = 0;
		rf_filter_coeff428_a = 0;
		rf_filter_coeff428_b = 0;
		rf_filter_coeff429_a = 0;
		rf_filter_coeff429_b = 0;
		rf_filter_coeff430_a = 0;
		rf_filter_coeff430_b = 0;
		rf_filter_coeff431_a = 0;
		rf_filter_coeff431_b = 0;
		rf_filter_coeff432_a = 0;
		rf_filter_coeff432_b = 0;
		rf_filter_coeff433_a = 0;
		rf_filter_coeff433_b = 0;
		rf_filter_coeff434_a = 0;
		rf_filter_coeff434_b = 0;
		rf_filter_coeff435_a = 0;
		rf_filter_coeff435_b = 0;
		rf_filter_coeff436_a = 0;
		rf_filter_coeff436_b = 0;
		rf_filter_coeff437_a = 0;
		rf_filter_coeff437_b = 0;
		rf_filter_coeff438_a = 0;
		rf_filter_coeff438_b = 0;
		rf_filter_coeff439_a = 0;
		rf_filter_coeff439_b = 0;
		rf_filter_coeff440_a = 0;
		rf_filter_coeff440_b = 0;
		rf_filter_coeff441_a = 0;
		rf_filter_coeff441_b = 0;
		rf_filter_coeff442_a = 0;
		rf_filter_coeff442_b = 0;
		rf_filter_coeff443_a = 0;
		rf_filter_coeff443_b = 0;
		rf_filter_coeff444_a = 0;
		rf_filter_coeff444_b = 0;
		rf_filter_coeff445_a = 0;
		rf_filter_coeff445_b = 0;
		rf_filter_coeff446_a = 0;
		rf_filter_coeff446_b = 0;
		rf_filter_coeff447_a = 0;
		rf_filter_coeff447_b = 0;
		rf_filter_coeff448_a = 0;
		rf_filter_coeff448_b = 0;
		rf_filter_coeff449_a = 0;
		rf_filter_coeff449_b = 0;
		rf_filter_coeff450_a = 0;
		rf_filter_coeff450_b = 0;
		rf_filter_coeff451_a = 0;
		rf_filter_coeff451_b = 0;
		rf_filter_coeff452_a = 0;
		rf_filter_coeff452_b = 0;
		rf_filter_coeff453_a = 0;
		rf_filter_coeff453_b = 0;
		rf_filter_coeff454_a = 0;
		rf_filter_coeff454_b = 0;
		rf_filter_coeff455_a = 0;
		rf_filter_coeff455_b = 0;
		rf_filter_coeff456_a = 0;
		rf_filter_coeff456_b = 0;
		rf_filter_coeff457_a = 0;
		rf_filter_coeff457_b = 0;
		rf_filter_coeff458_a = 0;
		rf_filter_coeff458_b = 0;
		rf_filter_coeff459_a = 0;
		rf_filter_coeff459_b = 0;
		rf_filter_coeff460_a = 0;
		rf_filter_coeff460_b = 0;
		rf_filter_coeff461_a = 0;
		rf_filter_coeff461_b = 0;
		rf_filter_coeff462_a = 0;
		rf_filter_coeff462_b = 0;
		rf_filter_coeff463_a = 0;
		rf_filter_coeff463_b = 0;
		rf_filter_coeff464_a = 0;
		rf_filter_coeff464_b = 0;
		rf_filter_coeff465_a = 0;
		rf_filter_coeff465_b = 0;
		rf_filter_coeff466_a = 0;
		rf_filter_coeff466_b = 0;
		rf_filter_coeff467_a = 0;
		rf_filter_coeff467_b = 0;
		rf_filter_coeff468_a = 0;
		rf_filter_coeff468_b = 0;
		rf_filter_coeff469_a = 0;
		rf_filter_coeff469_b = 0;
		rf_filter_coeff470_a = 0;
		rf_filter_coeff470_b = 0;
		rf_filter_coeff471_a = 0;
		rf_filter_coeff471_b = 0;
		rf_filter_coeff472_a = 0;
		rf_filter_coeff472_b = 0;
		rf_filter_coeff473_a = 0;
		rf_filter_coeff473_b = 0;
		rf_filter_coeff474_a = 0;
		rf_filter_coeff474_b = 0;
		rf_filter_coeff475_a = 0;
		rf_filter_coeff475_b = 0;
		rf_filter_coeff476_a = 0;
		rf_filter_coeff476_b = 0;
		rf_filter_coeff477_a = 0;
		rf_filter_coeff477_b = 0;
		rf_filter_coeff478_a = 0;
		rf_filter_coeff478_b = 0;
		rf_filter_coeff479_a = 0;
		rf_filter_coeff479_b = 0;
		rf_filter_coeff480_a = 0;
		rf_filter_coeff480_b = 0;
		rf_filter_coeff481_a = 0;
		rf_filter_coeff481_b = 0;
		rf_filter_coeff482_a = 0;
		rf_filter_coeff482_b = 0;
		rf_filter_coeff483_a = 0;
		rf_filter_coeff483_b = 0;
		rf_filter_coeff484_a = 0;
		rf_filter_coeff484_b = 0;
		rf_filter_coeff485_a = 0;
		rf_filter_coeff485_b = 0;
		rf_filter_coeff486_a = 0;
		rf_filter_coeff486_b = 0;
		rf_filter_coeff487_a = 0;
		rf_filter_coeff487_b = 0;
		rf_filter_coeff488_a = 0;
		rf_filter_coeff488_b = 0;
		rf_filter_coeff489_a = 0;
		rf_filter_coeff489_b = 0;
		rf_filter_coeff490_a = 0;
		rf_filter_coeff490_b = 0;
		rf_filter_coeff491_a = 0;
		rf_filter_coeff491_b = 0;
		rf_filter_coeff492_a = 0;
		rf_filter_coeff492_b = 0;
		rf_filter_coeff493_a = 0;
		rf_filter_coeff493_b = 0;
		rf_filter_coeff494_a = 0;
		rf_filter_coeff494_b = 0;
		rf_filter_coeff495_a = 0;
		rf_filter_coeff495_b = 0;
		rf_filter_coeff496_a = 0;
		rf_filter_coeff496_b = 0;
		rf_filter_coeff497_a = 0;
		rf_filter_coeff497_b = 0;
		rf_filter_coeff498_a = 0;
		rf_filter_coeff498_b = 0;
		rf_filter_coeff499_a = 0;
		rf_filter_coeff499_b = 0;
		rf_filter_coeff500_a = 0;
		rf_filter_coeff500_b = 0;
		rf_filter_coeff501_a = 0;
		rf_filter_coeff501_b = 0;
		rf_filter_coeff502_a = 0;
		rf_filter_coeff502_b = 0;
		rf_filter_coeff503_a = 0;
		rf_filter_coeff503_b = 0;
		rf_filter_coeff504_a = 0;
		rf_filter_coeff504_b = 0;
		rf_filter_coeff505_a = 0;
		rf_filter_coeff505_b = 0;
		rf_filter_coeff506_a = 0;
		rf_filter_coeff506_b = 0;
		rf_filter_coeff507_a = 0;
		rf_filter_coeff507_b = 0;
		rf_filter_coeff508_a = 0;
		rf_filter_coeff508_b = 0;
		rf_filter_coeff509_a = 0;
		rf_filter_coeff509_b = 0;
		rf_filter_coeff510_a = 0;
		rf_filter_coeff510_b = 0;
		rf_filter_coeff511_a = 0;
		rf_filter_coeff511_b = 0;

		// Wait 100 ns for global reset to finish
		#100;
		// Add stimulus here
		rstb = 1'b1;
		aud_in_rts = 1'b0;
		aud_out_rtr = 1'b0;
		#100;
		aud_in_rts = 1'b1;
		#5000;
		//aud_in_rts = 1'b0;
		#5000;
		aud_out_rtr = 1'b1;
		#100;
		//aud_out_rtr = 1'b0;
		filt_input_data = 32'hAAAAAAAA;
		
		
	end
	
	always
	begin
		forever #5 clk = ~clk;
	end
      
endmodule

