`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    13:04:49 06/06/2015 
// Design Name: 
// Module Name:    i2s_out 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module i2s_out(
    input clk,
    input rst,
    output sck,
    output ws,
    output sd,
    input [15:0] dout_lft,
    input [15:0] dout_rgt,
    input dout_rts,
    output dout_rtr,
    output fifo_overun
    );


endmodule
