//////////////////////////////////////////////////////////////////////////////////
// Module Name:             filter_mux.v
// Create Date:             ??? 
// Last Modification:       3/25/2016
// Author:                  Dhruvit Naik
// Description:             ????
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps
module filter_mux(clk, rden, rdptr, rddata,rf_filter_coeff0_a, rf_filter_coeff0_b,rf_filter_coeff1_a, rf_filter_coeff1_b,rf_filter_coeff2_a, rf_filter_coeff2_b,rf_filter_coeff3_a, rf_filter_coeff3_b,rf_filter_coeff4_a, rf_filter_coeff4_b,rf_filter_coeff5_a, rf_filter_coeff5_b,rf_filter_coeff6_a, rf_filter_coeff6_b,rf_filter_coeff7_a, rf_filter_coeff7_b,rf_filter_coeff8_a, rf_filter_coeff8_b,rf_filter_coeff9_a, rf_filter_coeff9_b,rf_filter_coeff10_a, rf_filter_coeff10_b,rf_filter_coeff11_a, rf_filter_coeff11_b,rf_filter_coeff12_a, rf_filter_coeff12_b,rf_filter_coeff13_a, rf_filter_coeff13_b,rf_filter_coeff14_a, rf_filter_coeff14_b,rf_filter_coeff15_a, rf_filter_coeff15_b,rf_filter_coeff16_a, rf_filter_coeff16_b,rf_filter_coeff17_a, rf_filter_coeff17_b,rf_filter_coeff18_a, rf_filter_coeff18_b,rf_filter_coeff19_a, rf_filter_coeff19_b,rf_filter_coeff20_a, rf_filter_coeff20_b,rf_filter_coeff21_a, rf_filter_coeff21_b,rf_filter_coeff22_a, rf_filter_coeff22_b,rf_filter_coeff23_a, rf_filter_coeff23_b,rf_filter_coeff24_a, rf_filter_coeff24_b,rf_filter_coeff25_a, rf_filter_coeff25_b,rf_filter_coeff26_a, rf_filter_coeff26_b,rf_filter_coeff27_a, rf_filter_coeff27_b,rf_filter_coeff28_a, rf_filter_coeff28_b,rf_filter_coeff29_a, rf_filter_coeff29_b,rf_filter_coeff30_a, rf_filter_coeff30_b,rf_filter_coeff31_a, rf_filter_coeff31_b,rf_filter_coeff32_a, rf_filter_coeff32_b,rf_filter_coeff33_a, rf_filter_coeff33_b,rf_filter_coeff34_a, rf_filter_coeff34_b,rf_filter_coeff35_a, rf_filter_coeff35_b,rf_filter_coeff36_a, rf_filter_coeff36_b,rf_filter_coeff37_a, rf_filter_coeff37_b,rf_filter_coeff38_a, rf_filter_coeff38_b,rf_filter_coeff39_a, rf_filter_coeff39_b,rf_filter_coeff40_a, rf_filter_coeff40_b,rf_filter_coeff41_a, rf_filter_coeff41_b,rf_filter_coeff42_a, rf_filter_coeff42_b,rf_filter_coeff43_a, rf_filter_coeff43_b,rf_filter_coeff44_a, rf_filter_coeff44_b,rf_filter_coeff45_a, rf_filter_coeff45_b,rf_filter_coeff46_a, rf_filter_coeff46_b,rf_filter_coeff47_a, rf_filter_coeff47_b,rf_filter_coeff48_a, rf_filter_coeff48_b,rf_filter_coeff49_a, rf_filter_coeff49_b,rf_filter_coeff50_a, rf_filter_coeff50_b,rf_filter_coeff51_a, rf_filter_coeff51_b,rf_filter_coeff52_a, rf_filter_coeff52_b,rf_filter_coeff53_a, rf_filter_coeff53_b,rf_filter_coeff54_a, rf_filter_coeff54_b,rf_filter_coeff55_a, rf_filter_coeff55_b,rf_filter_coeff56_a, rf_filter_coeff56_b,rf_filter_coeff57_a, rf_filter_coeff57_b,rf_filter_coeff58_a, rf_filter_coeff58_b,rf_filter_coeff59_a, rf_filter_coeff59_b,rf_filter_coeff60_a, rf_filter_coeff60_b,rf_filter_coeff61_a, rf_filter_coeff61_b,rf_filter_coeff62_a, rf_filter_coeff62_b,rf_filter_coeff63_a, rf_filter_coeff63_b,rf_filter_coeff64_a, rf_filter_coeff64_b,rf_filter_coeff65_a, rf_filter_coeff65_b,rf_filter_coeff66_a, rf_filter_coeff66_b,rf_filter_coeff67_a, rf_filter_coeff67_b,rf_filter_coeff68_a, rf_filter_coeff68_b,rf_filter_coeff69_a, rf_filter_coeff69_b,rf_filter_coeff70_a, rf_filter_coeff70_b,rf_filter_coeff71_a, rf_filter_coeff71_b,rf_filter_coeff72_a, rf_filter_coeff72_b,rf_filter_coeff73_a, rf_filter_coeff73_b,rf_filter_coeff74_a, rf_filter_coeff74_b,rf_filter_coeff75_a, rf_filter_coeff75_b,rf_filter_coeff76_a, rf_filter_coeff76_b,rf_filter_coeff77_a, rf_filter_coeff77_b,rf_filter_coeff78_a, rf_filter_coeff78_b,rf_filter_coeff79_a, rf_filter_coeff79_b,rf_filter_coeff80_a, rf_filter_coeff80_b,rf_filter_coeff81_a, rf_filter_coeff81_b,rf_filter_coeff82_a, rf_filter_coeff82_b,rf_filter_coeff83_a, rf_filter_coeff83_b,rf_filter_coeff84_a, rf_filter_coeff84_b,rf_filter_coeff85_a, rf_filter_coeff85_b,rf_filter_coeff86_a, rf_filter_coeff86_b,rf_filter_coeff87_a, rf_filter_coeff87_b,rf_filter_coeff88_a, rf_filter_coeff88_b,rf_filter_coeff89_a, rf_filter_coeff89_b,rf_filter_coeff90_a, rf_filter_coeff90_b,rf_filter_coeff91_a, rf_filter_coeff91_b,rf_filter_coeff92_a, rf_filter_coeff92_b,rf_filter_coeff93_a, rf_filter_coeff93_b,rf_filter_coeff94_a, rf_filter_coeff94_b,rf_filter_coeff95_a, rf_filter_coeff95_b,rf_filter_coeff96_a, rf_filter_coeff96_b,rf_filter_coeff97_a, rf_filter_coeff97_b,rf_filter_coeff98_a, rf_filter_coeff98_b,rf_filter_coeff99_a, rf_filter_coeff99_b,rf_filter_coeff100_a, rf_filter_coeff100_b,rf_filter_coeff101_a, rf_filter_coeff101_b,rf_filter_coeff102_a, rf_filter_coeff102_b,rf_filter_coeff103_a, rf_filter_coeff103_b,rf_filter_coeff104_a, rf_filter_coeff104_b,rf_filter_coeff105_a, rf_filter_coeff105_b,rf_filter_coeff106_a, rf_filter_coeff106_b,rf_filter_coeff107_a, rf_filter_coeff107_b,rf_filter_coeff108_a, rf_filter_coeff108_b,rf_filter_coeff109_a, rf_filter_coeff109_b,rf_filter_coeff110_a, rf_filter_coeff110_b,rf_filter_coeff111_a, rf_filter_coeff111_b,rf_filter_coeff112_a, rf_filter_coeff112_b,rf_filter_coeff113_a, rf_filter_coeff113_b,rf_filter_coeff114_a, rf_filter_coeff114_b,rf_filter_coeff115_a, rf_filter_coeff115_b,rf_filter_coeff116_a, rf_filter_coeff116_b,rf_filter_coeff117_a, rf_filter_coeff117_b,rf_filter_coeff118_a, rf_filter_coeff118_b,rf_filter_coeff119_a, rf_filter_coeff119_b,rf_filter_coeff120_a, rf_filter_coeff120_b,rf_filter_coeff121_a, rf_filter_coeff121_b,rf_filter_coeff122_a, rf_filter_coeff122_b,rf_filter_coeff123_a, rf_filter_coeff123_b,rf_filter_coeff124_a, rf_filter_coeff124_b,rf_filter_coeff125_a, rf_filter_coeff125_b,rf_filter_coeff126_a, rf_filter_coeff126_b,rf_filter_coeff127_a, rf_filter_coeff127_b,rf_filter_coeff128_a, rf_filter_coeff128_b,rf_filter_coeff129_a, rf_filter_coeff129_b,rf_filter_coeff130_a, rf_filter_coeff130_b,rf_filter_coeff131_a, rf_filter_coeff131_b,rf_filter_coeff132_a, rf_filter_coeff132_b,rf_filter_coeff133_a, rf_filter_coeff133_b,rf_filter_coeff134_a, rf_filter_coeff134_b,rf_filter_coeff135_a, rf_filter_coeff135_b,rf_filter_coeff136_a, rf_filter_coeff136_b,rf_filter_coeff137_a, rf_filter_coeff137_b,rf_filter_coeff138_a, rf_filter_coeff138_b,rf_filter_coeff139_a, rf_filter_coeff139_b,rf_filter_coeff140_a, rf_filter_coeff140_b,rf_filter_coeff141_a, rf_filter_coeff141_b,rf_filter_coeff142_a, rf_filter_coeff142_b,rf_filter_coeff143_a, rf_filter_coeff143_b,rf_filter_coeff144_a, rf_filter_coeff144_b,rf_filter_coeff145_a, rf_filter_coeff145_b,rf_filter_coeff146_a, rf_filter_coeff146_b,rf_filter_coeff147_a, rf_filter_coeff147_b,rf_filter_coeff148_a, rf_filter_coeff148_b,rf_filter_coeff149_a, rf_filter_coeff149_b,rf_filter_coeff150_a, rf_filter_coeff150_b,rf_filter_coeff151_a, rf_filter_coeff151_b,rf_filter_coeff152_a, rf_filter_coeff152_b,rf_filter_coeff153_a, rf_filter_coeff153_b,rf_filter_coeff154_a, rf_filter_coeff154_b,rf_filter_coeff155_a, rf_filter_coeff155_b,rf_filter_coeff156_a, rf_filter_coeff156_b,rf_filter_coeff157_a, rf_filter_coeff157_b,rf_filter_coeff158_a, rf_filter_coeff158_b,rf_filter_coeff159_a, rf_filter_coeff159_b,rf_filter_coeff160_a, rf_filter_coeff160_b,rf_filter_coeff161_a, rf_filter_coeff161_b,rf_filter_coeff162_a, rf_filter_coeff162_b,rf_filter_coeff163_a, rf_filter_coeff163_b,rf_filter_coeff164_a, rf_filter_coeff164_b,rf_filter_coeff165_a, rf_filter_coeff165_b,rf_filter_coeff166_a, rf_filter_coeff166_b,rf_filter_coeff167_a, rf_filter_coeff167_b,rf_filter_coeff168_a, rf_filter_coeff168_b,rf_filter_coeff169_a, rf_filter_coeff169_b,rf_filter_coeff170_a, rf_filter_coeff170_b,rf_filter_coeff171_a, rf_filter_coeff171_b,rf_filter_coeff172_a, rf_filter_coeff172_b,rf_filter_coeff173_a, rf_filter_coeff173_b,rf_filter_coeff174_a, rf_filter_coeff174_b,rf_filter_coeff175_a, rf_filter_coeff175_b,rf_filter_coeff176_a, rf_filter_coeff176_b,rf_filter_coeff177_a, rf_filter_coeff177_b,rf_filter_coeff178_a, rf_filter_coeff178_b,rf_filter_coeff179_a, rf_filter_coeff179_b,rf_filter_coeff180_a, rf_filter_coeff180_b,rf_filter_coeff181_a, rf_filter_coeff181_b,rf_filter_coeff182_a, rf_filter_coeff182_b,rf_filter_coeff183_a, rf_filter_coeff183_b,rf_filter_coeff184_a, rf_filter_coeff184_b,rf_filter_coeff185_a, rf_filter_coeff185_b,rf_filter_coeff186_a, rf_filter_coeff186_b,rf_filter_coeff187_a, rf_filter_coeff187_b,rf_filter_coeff188_a, rf_filter_coeff188_b,rf_filter_coeff189_a, rf_filter_coeff189_b,rf_filter_coeff190_a, rf_filter_coeff190_b,rf_filter_coeff191_a, rf_filter_coeff191_b,rf_filter_coeff192_a, rf_filter_coeff192_b,rf_filter_coeff193_a, rf_filter_coeff193_b,rf_filter_coeff194_a, rf_filter_coeff194_b,rf_filter_coeff195_a, rf_filter_coeff195_b,rf_filter_coeff196_a, rf_filter_coeff196_b,rf_filter_coeff197_a, rf_filter_coeff197_b,rf_filter_coeff198_a, rf_filter_coeff198_b,rf_filter_coeff199_a, rf_filter_coeff199_b,rf_filter_coeff200_a, rf_filter_coeff200_b,rf_filter_coeff201_a, rf_filter_coeff201_b,rf_filter_coeff202_a, rf_filter_coeff202_b,rf_filter_coeff203_a, rf_filter_coeff203_b,rf_filter_coeff204_a, rf_filter_coeff204_b,rf_filter_coeff205_a, rf_filter_coeff205_b,rf_filter_coeff206_a, rf_filter_coeff206_b,rf_filter_coeff207_a, rf_filter_coeff207_b,rf_filter_coeff208_a, rf_filter_coeff208_b,rf_filter_coeff209_a, rf_filter_coeff209_b,rf_filter_coeff210_a, rf_filter_coeff210_b,rf_filter_coeff211_a, rf_filter_coeff211_b,rf_filter_coeff212_a, rf_filter_coeff212_b,rf_filter_coeff213_a, rf_filter_coeff213_b,rf_filter_coeff214_a, rf_filter_coeff214_b,rf_filter_coeff215_a, rf_filter_coeff215_b,rf_filter_coeff216_a, rf_filter_coeff216_b,rf_filter_coeff217_a, rf_filter_coeff217_b,rf_filter_coeff218_a, rf_filter_coeff218_b,rf_filter_coeff219_a, rf_filter_coeff219_b,rf_filter_coeff220_a, rf_filter_coeff220_b,rf_filter_coeff221_a, rf_filter_coeff221_b,rf_filter_coeff222_a, rf_filter_coeff222_b,rf_filter_coeff223_a, rf_filter_coeff223_b,rf_filter_coeff224_a, rf_filter_coeff224_b,rf_filter_coeff225_a, rf_filter_coeff225_b,rf_filter_coeff226_a, rf_filter_coeff226_b,rf_filter_coeff227_a, rf_filter_coeff227_b,rf_filter_coeff228_a, rf_filter_coeff228_b,rf_filter_coeff229_a, rf_filter_coeff229_b,rf_filter_coeff230_a, rf_filter_coeff230_b,rf_filter_coeff231_a, rf_filter_coeff231_b,rf_filter_coeff232_a, rf_filter_coeff232_b,rf_filter_coeff233_a, rf_filter_coeff233_b,rf_filter_coeff234_a, rf_filter_coeff234_b,rf_filter_coeff235_a, rf_filter_coeff235_b,rf_filter_coeff236_a, rf_filter_coeff236_b,rf_filter_coeff237_a, rf_filter_coeff237_b,rf_filter_coeff238_a, rf_filter_coeff238_b,rf_filter_coeff239_a, rf_filter_coeff239_b,rf_filter_coeff240_a, rf_filter_coeff240_b,rf_filter_coeff241_a, rf_filter_coeff241_b,rf_filter_coeff242_a, rf_filter_coeff242_b,rf_filter_coeff243_a, rf_filter_coeff243_b,rf_filter_coeff244_a, rf_filter_coeff244_b,rf_filter_coeff245_a, rf_filter_coeff245_b,rf_filter_coeff246_a, rf_filter_coeff246_b,rf_filter_coeff247_a, rf_filter_coeff247_b,rf_filter_coeff248_a, rf_filter_coeff248_b,rf_filter_coeff249_a, rf_filter_coeff249_b,rf_filter_coeff250_a, rf_filter_coeff250_b,rf_filter_coeff251_a, rf_filter_coeff251_b,rf_filter_coeff252_a, rf_filter_coeff252_b,rf_filter_coeff253_a, rf_filter_coeff253_b,rf_filter_coeff254_a, rf_filter_coeff254_b,rf_filter_coeff255_a, rf_filter_coeff255_b,rf_filter_coeff256_a, rf_filter_coeff256_b,rf_filter_coeff257_a, rf_filter_coeff257_b,rf_filter_coeff258_a, rf_filter_coeff258_b,rf_filter_coeff259_a, rf_filter_coeff259_b,rf_filter_coeff260_a, rf_filter_coeff260_b,rf_filter_coeff261_a, rf_filter_coeff261_b,rf_filter_coeff262_a, rf_filter_coeff262_b,rf_filter_coeff263_a, rf_filter_coeff263_b,rf_filter_coeff264_a, rf_filter_coeff264_b,rf_filter_coeff265_a, rf_filter_coeff265_b,rf_filter_coeff266_a, rf_filter_coeff266_b,rf_filter_coeff267_a, rf_filter_coeff267_b,rf_filter_coeff268_a, rf_filter_coeff268_b,rf_filter_coeff269_a, rf_filter_coeff269_b,rf_filter_coeff270_a, rf_filter_coeff270_b,rf_filter_coeff271_a, rf_filter_coeff271_b,rf_filter_coeff272_a, rf_filter_coeff272_b,rf_filter_coeff273_a, rf_filter_coeff273_b,rf_filter_coeff274_a, rf_filter_coeff274_b,rf_filter_coeff275_a, rf_filter_coeff275_b,rf_filter_coeff276_a, rf_filter_coeff276_b,rf_filter_coeff277_a, rf_filter_coeff277_b,rf_filter_coeff278_a, rf_filter_coeff278_b,rf_filter_coeff279_a, rf_filter_coeff279_b,rf_filter_coeff280_a, rf_filter_coeff280_b,rf_filter_coeff281_a, rf_filter_coeff281_b,rf_filter_coeff282_a, rf_filter_coeff282_b,rf_filter_coeff283_a, rf_filter_coeff283_b,rf_filter_coeff284_a, rf_filter_coeff284_b,rf_filter_coeff285_a, rf_filter_coeff285_b,rf_filter_coeff286_a, rf_filter_coeff286_b,rf_filter_coeff287_a, rf_filter_coeff287_b,rf_filter_coeff288_a, rf_filter_coeff288_b,rf_filter_coeff289_a, rf_filter_coeff289_b,rf_filter_coeff290_a, rf_filter_coeff290_b,rf_filter_coeff291_a, rf_filter_coeff291_b,rf_filter_coeff292_a, rf_filter_coeff292_b,rf_filter_coeff293_a, rf_filter_coeff293_b,rf_filter_coeff294_a, rf_filter_coeff294_b,rf_filter_coeff295_a, rf_filter_coeff295_b,rf_filter_coeff296_a, rf_filter_coeff296_b,rf_filter_coeff297_a, rf_filter_coeff297_b,rf_filter_coeff298_a, rf_filter_coeff298_b,rf_filter_coeff299_a, rf_filter_coeff299_b,rf_filter_coeff300_a, rf_filter_coeff300_b,rf_filter_coeff301_a, rf_filter_coeff301_b,rf_filter_coeff302_a, rf_filter_coeff302_b,rf_filter_coeff303_a, rf_filter_coeff303_b,rf_filter_coeff304_a, rf_filter_coeff304_b,rf_filter_coeff305_a, rf_filter_coeff305_b,rf_filter_coeff306_a, rf_filter_coeff306_b,rf_filter_coeff307_a, rf_filter_coeff307_b,rf_filter_coeff308_a, rf_filter_coeff308_b,rf_filter_coeff309_a, rf_filter_coeff309_b,rf_filter_coeff310_a, rf_filter_coeff310_b,rf_filter_coeff311_a, rf_filter_coeff311_b,rf_filter_coeff312_a, rf_filter_coeff312_b,rf_filter_coeff313_a, rf_filter_coeff313_b,rf_filter_coeff314_a, rf_filter_coeff314_b,rf_filter_coeff315_a, rf_filter_coeff315_b,rf_filter_coeff316_a, rf_filter_coeff316_b,rf_filter_coeff317_a, rf_filter_coeff317_b,rf_filter_coeff318_a, rf_filter_coeff318_b,rf_filter_coeff319_a, rf_filter_coeff319_b,rf_filter_coeff320_a, rf_filter_coeff320_b,rf_filter_coeff321_a, rf_filter_coeff321_b,rf_filter_coeff322_a, rf_filter_coeff322_b,rf_filter_coeff323_a, rf_filter_coeff323_b,rf_filter_coeff324_a, rf_filter_coeff324_b,rf_filter_coeff325_a, rf_filter_coeff325_b,rf_filter_coeff326_a, rf_filter_coeff326_b,rf_filter_coeff327_a, rf_filter_coeff327_b,rf_filter_coeff328_a, rf_filter_coeff328_b,rf_filter_coeff329_a, rf_filter_coeff329_b,rf_filter_coeff330_a, rf_filter_coeff330_b,rf_filter_coeff331_a, rf_filter_coeff331_b,rf_filter_coeff332_a, rf_filter_coeff332_b,rf_filter_coeff333_a, rf_filter_coeff333_b,rf_filter_coeff334_a, rf_filter_coeff334_b,rf_filter_coeff335_a, rf_filter_coeff335_b,rf_filter_coeff336_a, rf_filter_coeff336_b,rf_filter_coeff337_a, rf_filter_coeff337_b,rf_filter_coeff338_a, rf_filter_coeff338_b,rf_filter_coeff339_a, rf_filter_coeff339_b,rf_filter_coeff340_a, rf_filter_coeff340_b,rf_filter_coeff341_a, rf_filter_coeff341_b,rf_filter_coeff342_a, rf_filter_coeff342_b,rf_filter_coeff343_a, rf_filter_coeff343_b,rf_filter_coeff344_a, rf_filter_coeff344_b,rf_filter_coeff345_a, rf_filter_coeff345_b,rf_filter_coeff346_a, rf_filter_coeff346_b,rf_filter_coeff347_a, rf_filter_coeff347_b,rf_filter_coeff348_a, rf_filter_coeff348_b,rf_filter_coeff349_a, rf_filter_coeff349_b,rf_filter_coeff350_a, rf_filter_coeff350_b,rf_filter_coeff351_a, rf_filter_coeff351_b,rf_filter_coeff352_a, rf_filter_coeff352_b,rf_filter_coeff353_a, rf_filter_coeff353_b,rf_filter_coeff354_a, rf_filter_coeff354_b,rf_filter_coeff355_a, rf_filter_coeff355_b,rf_filter_coeff356_a, rf_filter_coeff356_b,rf_filter_coeff357_a, rf_filter_coeff357_b,rf_filter_coeff358_a, rf_filter_coeff358_b,rf_filter_coeff359_a, rf_filter_coeff359_b,rf_filter_coeff360_a, rf_filter_coeff360_b,rf_filter_coeff361_a, rf_filter_coeff361_b,rf_filter_coeff362_a, rf_filter_coeff362_b,rf_filter_coeff363_a, rf_filter_coeff363_b,rf_filter_coeff364_a, rf_filter_coeff364_b,rf_filter_coeff365_a, rf_filter_coeff365_b,rf_filter_coeff366_a, rf_filter_coeff366_b,rf_filter_coeff367_a, rf_filter_coeff367_b,rf_filter_coeff368_a, rf_filter_coeff368_b,rf_filter_coeff369_a, rf_filter_coeff369_b,rf_filter_coeff370_a, rf_filter_coeff370_b,rf_filter_coeff371_a, rf_filter_coeff371_b,rf_filter_coeff372_a, rf_filter_coeff372_b,rf_filter_coeff373_a, rf_filter_coeff373_b,rf_filter_coeff374_a, rf_filter_coeff374_b,rf_filter_coeff375_a, rf_filter_coeff375_b,rf_filter_coeff376_a, rf_filter_coeff376_b,rf_filter_coeff377_a, rf_filter_coeff377_b,rf_filter_coeff378_a, rf_filter_coeff378_b,rf_filter_coeff379_a, rf_filter_coeff379_b,rf_filter_coeff380_a, rf_filter_coeff380_b,rf_filter_coeff381_a, rf_filter_coeff381_b,rf_filter_coeff382_a, rf_filter_coeff382_b,rf_filter_coeff383_a, rf_filter_coeff383_b,rf_filter_coeff384_a, rf_filter_coeff384_b,rf_filter_coeff385_a, rf_filter_coeff385_b,rf_filter_coeff386_a, rf_filter_coeff386_b,rf_filter_coeff387_a, rf_filter_coeff387_b,rf_filter_coeff388_a, rf_filter_coeff388_b,rf_filter_coeff389_a, rf_filter_coeff389_b,rf_filter_coeff390_a, rf_filter_coeff390_b,rf_filter_coeff391_a, rf_filter_coeff391_b,rf_filter_coeff392_a, rf_filter_coeff392_b,rf_filter_coeff393_a, rf_filter_coeff393_b,rf_filter_coeff394_a, rf_filter_coeff394_b,rf_filter_coeff395_a, rf_filter_coeff395_b,rf_filter_coeff396_a, rf_filter_coeff396_b,rf_filter_coeff397_a, rf_filter_coeff397_b,rf_filter_coeff398_a, rf_filter_coeff398_b,rf_filter_coeff399_a, rf_filter_coeff399_b,rf_filter_coeff400_a, rf_filter_coeff400_b,rf_filter_coeff401_a, rf_filter_coeff401_b,rf_filter_coeff402_a, rf_filter_coeff402_b,rf_filter_coeff403_a, rf_filter_coeff403_b,rf_filter_coeff404_a, rf_filter_coeff404_b,rf_filter_coeff405_a, rf_filter_coeff405_b,rf_filter_coeff406_a, rf_filter_coeff406_b,rf_filter_coeff407_a, rf_filter_coeff407_b,rf_filter_coeff408_a, rf_filter_coeff408_b,rf_filter_coeff409_a, rf_filter_coeff409_b,rf_filter_coeff410_a, rf_filter_coeff410_b,rf_filter_coeff411_a, rf_filter_coeff411_b,rf_filter_coeff412_a, rf_filter_coeff412_b,rf_filter_coeff413_a, rf_filter_coeff413_b,rf_filter_coeff414_a, rf_filter_coeff414_b,rf_filter_coeff415_a, rf_filter_coeff415_b,rf_filter_coeff416_a, rf_filter_coeff416_b,rf_filter_coeff417_a, rf_filter_coeff417_b,rf_filter_coeff418_a, rf_filter_coeff418_b,rf_filter_coeff419_a, rf_filter_coeff419_b,rf_filter_coeff420_a, rf_filter_coeff420_b,rf_filter_coeff421_a, rf_filter_coeff421_b,rf_filter_coeff422_a, rf_filter_coeff422_b,rf_filter_coeff423_a, rf_filter_coeff423_b,rf_filter_coeff424_a, rf_filter_coeff424_b,rf_filter_coeff425_a, rf_filter_coeff425_b,rf_filter_coeff426_a, rf_filter_coeff426_b,rf_filter_coeff427_a, rf_filter_coeff427_b,rf_filter_coeff428_a, rf_filter_coeff428_b,rf_filter_coeff429_a, rf_filter_coeff429_b,rf_filter_coeff430_a, rf_filter_coeff430_b,rf_filter_coeff431_a, rf_filter_coeff431_b,rf_filter_coeff432_a, rf_filter_coeff432_b,rf_filter_coeff433_a, rf_filter_coeff433_b,rf_filter_coeff434_a, rf_filter_coeff434_b,rf_filter_coeff435_a, rf_filter_coeff435_b,rf_filter_coeff436_a, rf_filter_coeff436_b,rf_filter_coeff437_a, rf_filter_coeff437_b,rf_filter_coeff438_a, rf_filter_coeff438_b,rf_filter_coeff439_a, rf_filter_coeff439_b,rf_filter_coeff440_a, rf_filter_coeff440_b,rf_filter_coeff441_a, rf_filter_coeff441_b,rf_filter_coeff442_a, rf_filter_coeff442_b,rf_filter_coeff443_a, rf_filter_coeff443_b,rf_filter_coeff444_a, rf_filter_coeff444_b,rf_filter_coeff445_a, rf_filter_coeff445_b,rf_filter_coeff446_a, rf_filter_coeff446_b,rf_filter_coeff447_a, rf_filter_coeff447_b,rf_filter_coeff448_a, rf_filter_coeff448_b,rf_filter_coeff449_a, rf_filter_coeff449_b,rf_filter_coeff450_a, rf_filter_coeff450_b,rf_filter_coeff451_a, rf_filter_coeff451_b,rf_filter_coeff452_a, rf_filter_coeff452_b,rf_filter_coeff453_a, rf_filter_coeff453_b,rf_filter_coeff454_a, rf_filter_coeff454_b,rf_filter_coeff455_a, rf_filter_coeff455_b,rf_filter_coeff456_a, rf_filter_coeff456_b,rf_filter_coeff457_a, rf_filter_coeff457_b,rf_filter_coeff458_a, rf_filter_coeff458_b,rf_filter_coeff459_a, rf_filter_coeff459_b,rf_filter_coeff460_a, rf_filter_coeff460_b,rf_filter_coeff461_a, rf_filter_coeff461_b,rf_filter_coeff462_a, rf_filter_coeff462_b,rf_filter_coeff463_a, rf_filter_coeff463_b,rf_filter_coeff464_a, rf_filter_coeff464_b,rf_filter_coeff465_a, rf_filter_coeff465_b,rf_filter_coeff466_a, rf_filter_coeff466_b,rf_filter_coeff467_a, rf_filter_coeff467_b,rf_filter_coeff468_a, rf_filter_coeff468_b,rf_filter_coeff469_a, rf_filter_coeff469_b,rf_filter_coeff470_a, rf_filter_coeff470_b,rf_filter_coeff471_a, rf_filter_coeff471_b,rf_filter_coeff472_a, rf_filter_coeff472_b,rf_filter_coeff473_a, rf_filter_coeff473_b,rf_filter_coeff474_a, rf_filter_coeff474_b,rf_filter_coeff475_a, rf_filter_coeff475_b,rf_filter_coeff476_a, rf_filter_coeff476_b,rf_filter_coeff477_a, rf_filter_coeff477_b,rf_filter_coeff478_a, rf_filter_coeff478_b,rf_filter_coeff479_a, rf_filter_coeff479_b,rf_filter_coeff480_a, rf_filter_coeff480_b,rf_filter_coeff481_a, rf_filter_coeff481_b,rf_filter_coeff482_a, rf_filter_coeff482_b,rf_filter_coeff483_a, rf_filter_coeff483_b,rf_filter_coeff484_a, rf_filter_coeff484_b,rf_filter_coeff485_a, rf_filter_coeff485_b,rf_filter_coeff486_a, rf_filter_coeff486_b,rf_filter_coeff487_a, rf_filter_coeff487_b,rf_filter_coeff488_a, rf_filter_coeff488_b,rf_filter_coeff489_a, rf_filter_coeff489_b,rf_filter_coeff490_a, rf_filter_coeff490_b,rf_filter_coeff491_a, rf_filter_coeff491_b,rf_filter_coeff492_a, rf_filter_coeff492_b,rf_filter_coeff493_a, rf_filter_coeff493_b,rf_filter_coeff494_a, rf_filter_coeff494_b,rf_filter_coeff495_a, rf_filter_coeff495_b,rf_filter_coeff496_a, rf_filter_coeff496_b,rf_filter_coeff497_a, rf_filter_coeff497_b,rf_filter_coeff498_a, rf_filter_coeff498_b,rf_filter_coeff499_a, rf_filter_coeff499_b,rf_filter_coeff500_a, rf_filter_coeff500_b,rf_filter_coeff501_a, rf_filter_coeff501_b,rf_filter_coeff502_a, rf_filter_coeff502_b,rf_filter_coeff503_a, rf_filter_coeff503_b,rf_filter_coeff504_a, rf_filter_coeff504_b,rf_filter_coeff505_a, rf_filter_coeff505_b,rf_filter_coeff506_a, rf_filter_coeff506_b,rf_filter_coeff507_a, rf_filter_coeff507_b,rf_filter_coeff508_a, rf_filter_coeff508_b,rf_filter_coeff509_a, rf_filter_coeff509_b,rf_filter_coeff510_a, rf_filter_coeff510_b,rf_filter_coeff511_a, rf_filter_coeff511_b
   );

    input [7:0] rf_filter_coeff0_a, rf_filter_coeff0_b,
    rf_filter_coeff1_a, rf_filter_coeff1_b,rf_filter_coeff2_a, rf_filter_coeff2_b,rf_filter_coeff3_a, rf_filter_coeff3_b,rf_filter_coeff4_a, rf_filter_coeff4_b,
    rf_filter_coeff5_a, rf_filter_coeff5_b,rf_filter_coeff6_a, rf_filter_coeff6_b,rf_filter_coeff7_a, rf_filter_coeff7_b,rf_filter_coeff8_a, rf_filter_coeff8_b,
    rf_filter_coeff9_a, rf_filter_coeff9_b,rf_filter_coeff10_a, rf_filter_coeff10_b,rf_filter_coeff11_a, rf_filter_coeff11_b,rf_filter_coeff12_a, rf_filter_coeff12_b,
    rf_filter_coeff13_a, rf_filter_coeff13_b,rf_filter_coeff14_a, rf_filter_coeff14_b,rf_filter_coeff15_a, rf_filter_coeff15_b,rf_filter_coeff16_a, rf_filter_coeff16_b,
    rf_filter_coeff17_a, rf_filter_coeff17_b,rf_filter_coeff18_a, rf_filter_coeff18_b,rf_filter_coeff19_a, rf_filter_coeff19_b,rf_filter_coeff20_a, rf_filter_coeff20_b,
    rf_filter_coeff21_a, rf_filter_coeff21_b,rf_filter_coeff22_a, rf_filter_coeff22_b,rf_filter_coeff23_a, rf_filter_coeff23_b,rf_filter_coeff24_a, rf_filter_coeff24_b,
    rf_filter_coeff25_a, rf_filter_coeff25_b,rf_filter_coeff26_a, rf_filter_coeff26_b,rf_filter_coeff27_a, rf_filter_coeff27_b,rf_filter_coeff28_a, rf_filter_coeff28_b,
    rf_filter_coeff29_a, rf_filter_coeff29_b,rf_filter_coeff30_a, rf_filter_coeff30_b,rf_filter_coeff31_a, rf_filter_coeff31_b,rf_filter_coeff32_a, rf_filter_coeff32_b,
    rf_filter_coeff33_a, rf_filter_coeff33_b,rf_filter_coeff34_a, rf_filter_coeff34_b,rf_filter_coeff35_a, rf_filter_coeff35_b,rf_filter_coeff36_a, rf_filter_coeff36_b,
    rf_filter_coeff37_a, rf_filter_coeff37_b,rf_filter_coeff38_a, rf_filter_coeff38_b,rf_filter_coeff39_a, rf_filter_coeff39_b,rf_filter_coeff40_a, rf_filter_coeff40_b,
    rf_filter_coeff41_a, rf_filter_coeff41_b,rf_filter_coeff42_a, rf_filter_coeff42_b,rf_filter_coeff43_a, rf_filter_coeff43_b,rf_filter_coeff44_a, rf_filter_coeff44_b,
    rf_filter_coeff45_a, rf_filter_coeff45_b,rf_filter_coeff46_a, rf_filter_coeff46_b,rf_filter_coeff47_a, rf_filter_coeff47_b,rf_filter_coeff48_a, rf_filter_coeff48_b,
    rf_filter_coeff49_a, rf_filter_coeff49_b,rf_filter_coeff50_a, rf_filter_coeff50_b,rf_filter_coeff51_a, rf_filter_coeff51_b,rf_filter_coeff52_a, rf_filter_coeff52_b,
    rf_filter_coeff53_a, rf_filter_coeff53_b,rf_filter_coeff54_a, rf_filter_coeff54_b,rf_filter_coeff55_a, rf_filter_coeff55_b,rf_filter_coeff56_a, rf_filter_coeff56_b,
    rf_filter_coeff57_a, rf_filter_coeff57_b,rf_filter_coeff58_a, rf_filter_coeff58_b,rf_filter_coeff59_a, rf_filter_coeff59_b,rf_filter_coeff60_a, rf_filter_coeff60_b,
    rf_filter_coeff61_a, rf_filter_coeff61_b,rf_filter_coeff62_a, rf_filter_coeff62_b,rf_filter_coeff63_a, rf_filter_coeff63_b,rf_filter_coeff64_a, rf_filter_coeff64_b,
    rf_filter_coeff65_a, rf_filter_coeff65_b,rf_filter_coeff66_a, rf_filter_coeff66_b,rf_filter_coeff67_a, rf_filter_coeff67_b,rf_filter_coeff68_a, rf_filter_coeff68_b,
    rf_filter_coeff69_a, rf_filter_coeff69_b,rf_filter_coeff70_a, rf_filter_coeff70_b,rf_filter_coeff71_a, rf_filter_coeff71_b,rf_filter_coeff72_a, rf_filter_coeff72_b,
    rf_filter_coeff73_a, rf_filter_coeff73_b,rf_filter_coeff74_a, rf_filter_coeff74_b,rf_filter_coeff75_a, rf_filter_coeff75_b,rf_filter_coeff76_a, rf_filter_coeff76_b,
    rf_filter_coeff77_a, rf_filter_coeff77_b,rf_filter_coeff78_a, rf_filter_coeff78_b,rf_filter_coeff79_a, rf_filter_coeff79_b,rf_filter_coeff80_a, rf_filter_coeff80_b,
    rf_filter_coeff81_a, rf_filter_coeff81_b,rf_filter_coeff82_a, rf_filter_coeff82_b,rf_filter_coeff83_a, rf_filter_coeff83_b,rf_filter_coeff84_a, rf_filter_coeff84_b,
    rf_filter_coeff85_a, rf_filter_coeff85_b,rf_filter_coeff86_a, rf_filter_coeff86_b,rf_filter_coeff87_a, rf_filter_coeff87_b,rf_filter_coeff88_a, rf_filter_coeff88_b,
    rf_filter_coeff89_a, rf_filter_coeff89_b,rf_filter_coeff90_a, rf_filter_coeff90_b,rf_filter_coeff91_a, rf_filter_coeff91_b,rf_filter_coeff92_a, rf_filter_coeff92_b,
    rf_filter_coeff93_a, rf_filter_coeff93_b,rf_filter_coeff94_a, rf_filter_coeff94_b,rf_filter_coeff95_a, rf_filter_coeff95_b,rf_filter_coeff96_a, rf_filter_coeff96_b,
    rf_filter_coeff97_a, rf_filter_coeff97_b,rf_filter_coeff98_a, rf_filter_coeff98_b,rf_filter_coeff99_a, rf_filter_coeff99_b,rf_filter_coeff100_a, rf_filter_coeff100_b,
    rf_filter_coeff101_a, rf_filter_coeff101_b,rf_filter_coeff102_a, rf_filter_coeff102_b,rf_filter_coeff103_a, rf_filter_coeff103_b,rf_filter_coeff104_a, rf_filter_coeff104_b,
    rf_filter_coeff105_a, rf_filter_coeff105_b,rf_filter_coeff106_a, rf_filter_coeff106_b,rf_filter_coeff107_a, rf_filter_coeff107_b,rf_filter_coeff108_a, rf_filter_coeff108_b,
    rf_filter_coeff109_a, rf_filter_coeff109_b,rf_filter_coeff110_a, rf_filter_coeff110_b,rf_filter_coeff111_a, rf_filter_coeff111_b,rf_filter_coeff112_a, rf_filter_coeff112_b,
    rf_filter_coeff113_a, rf_filter_coeff113_b,rf_filter_coeff114_a, rf_filter_coeff114_b,rf_filter_coeff115_a, rf_filter_coeff115_b,rf_filter_coeff116_a, rf_filter_coeff116_b,
    rf_filter_coeff117_a, rf_filter_coeff117_b,rf_filter_coeff118_a, rf_filter_coeff118_b,rf_filter_coeff119_a, rf_filter_coeff119_b,rf_filter_coeff120_a, rf_filter_coeff120_b,
    rf_filter_coeff121_a, rf_filter_coeff121_b,rf_filter_coeff122_a, rf_filter_coeff122_b,rf_filter_coeff123_a, rf_filter_coeff123_b,rf_filter_coeff124_a, rf_filter_coeff124_b,
    rf_filter_coeff125_a, rf_filter_coeff125_b,rf_filter_coeff126_a, rf_filter_coeff126_b,rf_filter_coeff127_a, rf_filter_coeff127_b,rf_filter_coeff128_a, rf_filter_coeff128_b,
    rf_filter_coeff129_a, rf_filter_coeff129_b,rf_filter_coeff130_a, rf_filter_coeff130_b,rf_filter_coeff131_a, rf_filter_coeff131_b,rf_filter_coeff132_a, rf_filter_coeff132_b,
    rf_filter_coeff133_a, rf_filter_coeff133_b,rf_filter_coeff134_a, rf_filter_coeff134_b,rf_filter_coeff135_a, rf_filter_coeff135_b,rf_filter_coeff136_a, rf_filter_coeff136_b,
    rf_filter_coeff137_a, rf_filter_coeff137_b,rf_filter_coeff138_a, rf_filter_coeff138_b,rf_filter_coeff139_a, rf_filter_coeff139_b,rf_filter_coeff140_a, rf_filter_coeff140_b,
    rf_filter_coeff141_a, rf_filter_coeff141_b,rf_filter_coeff142_a, rf_filter_coeff142_b,rf_filter_coeff143_a, rf_filter_coeff143_b,rf_filter_coeff144_a, rf_filter_coeff144_b,
    rf_filter_coeff145_a, rf_filter_coeff145_b,rf_filter_coeff146_a, rf_filter_coeff146_b,rf_filter_coeff147_a, rf_filter_coeff147_b,rf_filter_coeff148_a, rf_filter_coeff148_b,
    rf_filter_coeff149_a, rf_filter_coeff149_b,rf_filter_coeff150_a, rf_filter_coeff150_b,rf_filter_coeff151_a, rf_filter_coeff151_b,rf_filter_coeff152_a, rf_filter_coeff152_b,
    rf_filter_coeff153_a, rf_filter_coeff153_b,rf_filter_coeff154_a, rf_filter_coeff154_b,rf_filter_coeff155_a, rf_filter_coeff155_b,rf_filter_coeff156_a, rf_filter_coeff156_b,
    rf_filter_coeff157_a, rf_filter_coeff157_b,rf_filter_coeff158_a, rf_filter_coeff158_b,rf_filter_coeff159_a, rf_filter_coeff159_b,rf_filter_coeff160_a, rf_filter_coeff160_b,
    rf_filter_coeff161_a, rf_filter_coeff161_b,rf_filter_coeff162_a, rf_filter_coeff162_b,rf_filter_coeff163_a, rf_filter_coeff163_b,rf_filter_coeff164_a, rf_filter_coeff164_b,
    rf_filter_coeff165_a, rf_filter_coeff165_b,rf_filter_coeff166_a, rf_filter_coeff166_b,rf_filter_coeff167_a, rf_filter_coeff167_b,rf_filter_coeff168_a, rf_filter_coeff168_b,
    rf_filter_coeff169_a, rf_filter_coeff169_b,rf_filter_coeff170_a, rf_filter_coeff170_b,rf_filter_coeff171_a, rf_filter_coeff171_b,rf_filter_coeff172_a, rf_filter_coeff172_b,
    rf_filter_coeff173_a, rf_filter_coeff173_b,rf_filter_coeff174_a, rf_filter_coeff174_b,rf_filter_coeff175_a, rf_filter_coeff175_b,rf_filter_coeff176_a, rf_filter_coeff176_b,
    rf_filter_coeff177_a, rf_filter_coeff177_b,rf_filter_coeff178_a, rf_filter_coeff178_b,rf_filter_coeff179_a, rf_filter_coeff179_b,rf_filter_coeff180_a, rf_filter_coeff180_b,
    rf_filter_coeff181_a, rf_filter_coeff181_b,rf_filter_coeff182_a, rf_filter_coeff182_b,rf_filter_coeff183_a, rf_filter_coeff183_b,rf_filter_coeff184_a, rf_filter_coeff184_b,
    rf_filter_coeff185_a, rf_filter_coeff185_b,rf_filter_coeff186_a, rf_filter_coeff186_b,rf_filter_coeff187_a, rf_filter_coeff187_b,rf_filter_coeff188_a, rf_filter_coeff188_b,
    rf_filter_coeff189_a, rf_filter_coeff189_b,rf_filter_coeff190_a, rf_filter_coeff190_b,rf_filter_coeff191_a, rf_filter_coeff191_b,rf_filter_coeff192_a, rf_filter_coeff192_b,
    rf_filter_coeff193_a, rf_filter_coeff193_b,rf_filter_coeff194_a, rf_filter_coeff194_b,rf_filter_coeff195_a, rf_filter_coeff195_b,rf_filter_coeff196_a, rf_filter_coeff196_b,
    rf_filter_coeff197_a, rf_filter_coeff197_b,rf_filter_coeff198_a, rf_filter_coeff198_b,rf_filter_coeff199_a, rf_filter_coeff199_b,rf_filter_coeff200_a, rf_filter_coeff200_b,
    rf_filter_coeff201_a, rf_filter_coeff201_b,rf_filter_coeff202_a, rf_filter_coeff202_b,rf_filter_coeff203_a, rf_filter_coeff203_b,rf_filter_coeff204_a, rf_filter_coeff204_b,
    rf_filter_coeff205_a, rf_filter_coeff205_b,rf_filter_coeff206_a, rf_filter_coeff206_b,rf_filter_coeff207_a, rf_filter_coeff207_b,rf_filter_coeff208_a, rf_filter_coeff208_b,
    rf_filter_coeff209_a, rf_filter_coeff209_b,rf_filter_coeff210_a, rf_filter_coeff210_b,rf_filter_coeff211_a, rf_filter_coeff211_b,rf_filter_coeff212_a, rf_filter_coeff212_b,
    rf_filter_coeff213_a, rf_filter_coeff213_b,rf_filter_coeff214_a, rf_filter_coeff214_b,rf_filter_coeff215_a, rf_filter_coeff215_b,rf_filter_coeff216_a, rf_filter_coeff216_b,
    rf_filter_coeff217_a, rf_filter_coeff217_b,rf_filter_coeff218_a, rf_filter_coeff218_b,rf_filter_coeff219_a, rf_filter_coeff219_b,rf_filter_coeff220_a, rf_filter_coeff220_b,
    rf_filter_coeff221_a, rf_filter_coeff221_b,rf_filter_coeff222_a, rf_filter_coeff222_b,rf_filter_coeff223_a, rf_filter_coeff223_b,rf_filter_coeff224_a, rf_filter_coeff224_b,
    rf_filter_coeff225_a, rf_filter_coeff225_b,rf_filter_coeff226_a, rf_filter_coeff226_b,rf_filter_coeff227_a, rf_filter_coeff227_b,rf_filter_coeff228_a, rf_filter_coeff228_b,
    rf_filter_coeff229_a, rf_filter_coeff229_b,rf_filter_coeff230_a, rf_filter_coeff230_b,rf_filter_coeff231_a, rf_filter_coeff231_b,rf_filter_coeff232_a, rf_filter_coeff232_b,
    rf_filter_coeff233_a, rf_filter_coeff233_b,rf_filter_coeff234_a, rf_filter_coeff234_b,rf_filter_coeff235_a, rf_filter_coeff235_b,rf_filter_coeff236_a, rf_filter_coeff236_b,
    rf_filter_coeff237_a, rf_filter_coeff237_b,rf_filter_coeff238_a, rf_filter_coeff238_b,rf_filter_coeff239_a, rf_filter_coeff239_b,rf_filter_coeff240_a, rf_filter_coeff240_b,
    rf_filter_coeff241_a, rf_filter_coeff241_b,rf_filter_coeff242_a, rf_filter_coeff242_b,rf_filter_coeff243_a, rf_filter_coeff243_b,rf_filter_coeff244_a, rf_filter_coeff244_b,
    rf_filter_coeff245_a, rf_filter_coeff245_b,rf_filter_coeff246_a, rf_filter_coeff246_b,rf_filter_coeff247_a, rf_filter_coeff247_b,rf_filter_coeff248_a, rf_filter_coeff248_b,
    rf_filter_coeff249_a, rf_filter_coeff249_b,rf_filter_coeff250_a, rf_filter_coeff250_b,rf_filter_coeff251_a, rf_filter_coeff251_b,rf_filter_coeff252_a, rf_filter_coeff252_b,
    rf_filter_coeff253_a, rf_filter_coeff253_b,rf_filter_coeff254_a, rf_filter_coeff254_b,rf_filter_coeff255_a, rf_filter_coeff255_b,rf_filter_coeff256_a, rf_filter_coeff256_b,
    rf_filter_coeff257_a, rf_filter_coeff257_b,rf_filter_coeff258_a, rf_filter_coeff258_b,rf_filter_coeff259_a, rf_filter_coeff259_b,rf_filter_coeff260_a, rf_filter_coeff260_b,
    rf_filter_coeff261_a, rf_filter_coeff261_b,rf_filter_coeff262_a, rf_filter_coeff262_b,rf_filter_coeff263_a, rf_filter_coeff263_b,rf_filter_coeff264_a, rf_filter_coeff264_b,
    rf_filter_coeff265_a, rf_filter_coeff265_b,rf_filter_coeff266_a, rf_filter_coeff266_b,rf_filter_coeff267_a, rf_filter_coeff267_b,rf_filter_coeff268_a, rf_filter_coeff268_b,
    rf_filter_coeff269_a, rf_filter_coeff269_b,rf_filter_coeff270_a, rf_filter_coeff270_b,rf_filter_coeff271_a, rf_filter_coeff271_b,rf_filter_coeff272_a, rf_filter_coeff272_b,
    rf_filter_coeff273_a, rf_filter_coeff273_b,rf_filter_coeff274_a, rf_filter_coeff274_b,rf_filter_coeff275_a, rf_filter_coeff275_b,rf_filter_coeff276_a, rf_filter_coeff276_b,
    rf_filter_coeff277_a, rf_filter_coeff277_b,rf_filter_coeff278_a, rf_filter_coeff278_b,rf_filter_coeff279_a, rf_filter_coeff279_b,rf_filter_coeff280_a, rf_filter_coeff280_b,
    rf_filter_coeff281_a, rf_filter_coeff281_b,rf_filter_coeff282_a, rf_filter_coeff282_b,rf_filter_coeff283_a, rf_filter_coeff283_b,rf_filter_coeff284_a, rf_filter_coeff284_b,
    rf_filter_coeff285_a, rf_filter_coeff285_b,rf_filter_coeff286_a, rf_filter_coeff286_b,rf_filter_coeff287_a, rf_filter_coeff287_b,rf_filter_coeff288_a, rf_filter_coeff288_b,
    rf_filter_coeff289_a, rf_filter_coeff289_b,rf_filter_coeff290_a, rf_filter_coeff290_b,rf_filter_coeff291_a, rf_filter_coeff291_b,rf_filter_coeff292_a, rf_filter_coeff292_b,
    rf_filter_coeff293_a, rf_filter_coeff293_b,rf_filter_coeff294_a, rf_filter_coeff294_b,rf_filter_coeff295_a, rf_filter_coeff295_b,rf_filter_coeff296_a, rf_filter_coeff296_b,
    rf_filter_coeff297_a, rf_filter_coeff297_b,rf_filter_coeff298_a, rf_filter_coeff298_b,rf_filter_coeff299_a, rf_filter_coeff299_b,rf_filter_coeff300_a, rf_filter_coeff300_b,
    rf_filter_coeff301_a, rf_filter_coeff301_b,rf_filter_coeff302_a, rf_filter_coeff302_b,rf_filter_coeff303_a, rf_filter_coeff303_b,rf_filter_coeff304_a, rf_filter_coeff304_b,
    rf_filter_coeff305_a, rf_filter_coeff305_b,rf_filter_coeff306_a, rf_filter_coeff306_b,rf_filter_coeff307_a, rf_filter_coeff307_b,rf_filter_coeff308_a, rf_filter_coeff308_b,
    rf_filter_coeff309_a, rf_filter_coeff309_b,rf_filter_coeff310_a, rf_filter_coeff310_b,rf_filter_coeff311_a, rf_filter_coeff311_b,rf_filter_coeff312_a, rf_filter_coeff312_b,
    rf_filter_coeff313_a, rf_filter_coeff313_b,rf_filter_coeff314_a, rf_filter_coeff314_b,rf_filter_coeff315_a, rf_filter_coeff315_b,rf_filter_coeff316_a, rf_filter_coeff316_b,
    rf_filter_coeff317_a, rf_filter_coeff317_b,rf_filter_coeff318_a, rf_filter_coeff318_b,rf_filter_coeff319_a, rf_filter_coeff319_b,rf_filter_coeff320_a, rf_filter_coeff320_b,
    rf_filter_coeff321_a, rf_filter_coeff321_b,rf_filter_coeff322_a, rf_filter_coeff322_b,rf_filter_coeff323_a, rf_filter_coeff323_b,rf_filter_coeff324_a, rf_filter_coeff324_b,
    rf_filter_coeff325_a, rf_filter_coeff325_b,rf_filter_coeff326_a, rf_filter_coeff326_b,rf_filter_coeff327_a, rf_filter_coeff327_b,rf_filter_coeff328_a, rf_filter_coeff328_b,
    rf_filter_coeff329_a, rf_filter_coeff329_b,rf_filter_coeff330_a, rf_filter_coeff330_b,rf_filter_coeff331_a, rf_filter_coeff331_b,rf_filter_coeff332_a, rf_filter_coeff332_b,
    rf_filter_coeff333_a, rf_filter_coeff333_b,rf_filter_coeff334_a, rf_filter_coeff334_b,rf_filter_coeff335_a, rf_filter_coeff335_b,rf_filter_coeff336_a, rf_filter_coeff336_b,
    rf_filter_coeff337_a, rf_filter_coeff337_b,rf_filter_coeff338_a, rf_filter_coeff338_b,rf_filter_coeff339_a, rf_filter_coeff339_b,rf_filter_coeff340_a, rf_filter_coeff340_b,
    rf_filter_coeff341_a, rf_filter_coeff341_b,rf_filter_coeff342_a, rf_filter_coeff342_b,rf_filter_coeff343_a, rf_filter_coeff343_b,rf_filter_coeff344_a, rf_filter_coeff344_b,
    rf_filter_coeff345_a, rf_filter_coeff345_b,rf_filter_coeff346_a, rf_filter_coeff346_b,rf_filter_coeff347_a, rf_filter_coeff347_b,rf_filter_coeff348_a, rf_filter_coeff348_b,
    rf_filter_coeff349_a, rf_filter_coeff349_b,rf_filter_coeff350_a, rf_filter_coeff350_b,rf_filter_coeff351_a, rf_filter_coeff351_b,rf_filter_coeff352_a, rf_filter_coeff352_b,
    rf_filter_coeff353_a, rf_filter_coeff353_b,rf_filter_coeff354_a, rf_filter_coeff354_b,rf_filter_coeff355_a, rf_filter_coeff355_b,rf_filter_coeff356_a, rf_filter_coeff356_b,
    rf_filter_coeff357_a, rf_filter_coeff357_b,rf_filter_coeff358_a, rf_filter_coeff358_b,rf_filter_coeff359_a, rf_filter_coeff359_b,rf_filter_coeff360_a, rf_filter_coeff360_b,
    rf_filter_coeff361_a, rf_filter_coeff361_b,rf_filter_coeff362_a, rf_filter_coeff362_b,rf_filter_coeff363_a, rf_filter_coeff363_b,rf_filter_coeff364_a, rf_filter_coeff364_b,
    rf_filter_coeff365_a, rf_filter_coeff365_b,rf_filter_coeff366_a, rf_filter_coeff366_b,rf_filter_coeff367_a, rf_filter_coeff367_b,rf_filter_coeff368_a, rf_filter_coeff368_b,
    rf_filter_coeff369_a, rf_filter_coeff369_b,rf_filter_coeff370_a, rf_filter_coeff370_b,rf_filter_coeff371_a, rf_filter_coeff371_b,rf_filter_coeff372_a, rf_filter_coeff372_b,
    rf_filter_coeff373_a, rf_filter_coeff373_b,rf_filter_coeff374_a, rf_filter_coeff374_b,rf_filter_coeff375_a, rf_filter_coeff375_b,rf_filter_coeff376_a, rf_filter_coeff376_b,
    rf_filter_coeff377_a, rf_filter_coeff377_b,rf_filter_coeff378_a, rf_filter_coeff378_b,rf_filter_coeff379_a, rf_filter_coeff379_b,rf_filter_coeff380_a, rf_filter_coeff380_b,
    rf_filter_coeff381_a, rf_filter_coeff381_b,rf_filter_coeff382_a, rf_filter_coeff382_b,rf_filter_coeff383_a, rf_filter_coeff383_b,rf_filter_coeff384_a, rf_filter_coeff384_b,
    rf_filter_coeff385_a, rf_filter_coeff385_b,rf_filter_coeff386_a, rf_filter_coeff386_b,rf_filter_coeff387_a, rf_filter_coeff387_b,rf_filter_coeff388_a, rf_filter_coeff388_b,
    rf_filter_coeff389_a, rf_filter_coeff389_b,rf_filter_coeff390_a, rf_filter_coeff390_b,rf_filter_coeff391_a, rf_filter_coeff391_b,rf_filter_coeff392_a, rf_filter_coeff392_b,
    rf_filter_coeff393_a, rf_filter_coeff393_b,rf_filter_coeff394_a, rf_filter_coeff394_b,rf_filter_coeff395_a, rf_filter_coeff395_b,rf_filter_coeff396_a, rf_filter_coeff396_b,
    rf_filter_coeff397_a, rf_filter_coeff397_b,rf_filter_coeff398_a, rf_filter_coeff398_b,rf_filter_coeff399_a, rf_filter_coeff399_b,rf_filter_coeff400_a, rf_filter_coeff400_b,
    rf_filter_coeff401_a, rf_filter_coeff401_b,rf_filter_coeff402_a, rf_filter_coeff402_b,rf_filter_coeff403_a, rf_filter_coeff403_b,rf_filter_coeff404_a, rf_filter_coeff404_b,
    rf_filter_coeff405_a, rf_filter_coeff405_b,rf_filter_coeff406_a, rf_filter_coeff406_b,rf_filter_coeff407_a, rf_filter_coeff407_b,rf_filter_coeff408_a, rf_filter_coeff408_b,
    rf_filter_coeff409_a, rf_filter_coeff409_b,rf_filter_coeff410_a, rf_filter_coeff410_b,rf_filter_coeff411_a, rf_filter_coeff411_b,rf_filter_coeff412_a, rf_filter_coeff412_b,
    rf_filter_coeff413_a, rf_filter_coeff413_b,rf_filter_coeff414_a, rf_filter_coeff414_b,rf_filter_coeff415_a, rf_filter_coeff415_b,rf_filter_coeff416_a, rf_filter_coeff416_b,
    rf_filter_coeff417_a, rf_filter_coeff417_b,rf_filter_coeff418_a, rf_filter_coeff418_b,rf_filter_coeff419_a, rf_filter_coeff419_b,rf_filter_coeff420_a, rf_filter_coeff420_b,
    rf_filter_coeff421_a, rf_filter_coeff421_b,rf_filter_coeff422_a, rf_filter_coeff422_b,rf_filter_coeff423_a, rf_filter_coeff423_b,rf_filter_coeff424_a, rf_filter_coeff424_b,
    rf_filter_coeff425_a, rf_filter_coeff425_b,rf_filter_coeff426_a, rf_filter_coeff426_b,rf_filter_coeff427_a, rf_filter_coeff427_b,rf_filter_coeff428_a, rf_filter_coeff428_b,
    rf_filter_coeff429_a, rf_filter_coeff429_b,rf_filter_coeff430_a, rf_filter_coeff430_b,rf_filter_coeff431_a, rf_filter_coeff431_b,rf_filter_coeff432_a, rf_filter_coeff432_b,
    rf_filter_coeff433_a, rf_filter_coeff433_b,rf_filter_coeff434_a, rf_filter_coeff434_b,rf_filter_coeff435_a, rf_filter_coeff435_b,rf_filter_coeff436_a, rf_filter_coeff436_b,
    rf_filter_coeff437_a, rf_filter_coeff437_b,rf_filter_coeff438_a, rf_filter_coeff438_b,rf_filter_coeff439_a, rf_filter_coeff439_b,rf_filter_coeff440_a, rf_filter_coeff440_b,
    rf_filter_coeff441_a, rf_filter_coeff441_b,rf_filter_coeff442_a, rf_filter_coeff442_b,rf_filter_coeff443_a, rf_filter_coeff443_b,rf_filter_coeff444_a, rf_filter_coeff444_b,
    rf_filter_coeff445_a, rf_filter_coeff445_b,rf_filter_coeff446_a, rf_filter_coeff446_b,rf_filter_coeff447_a, rf_filter_coeff447_b,rf_filter_coeff448_a, rf_filter_coeff448_b,
    rf_filter_coeff449_a, rf_filter_coeff449_b,rf_filter_coeff450_a, rf_filter_coeff450_b,rf_filter_coeff451_a, rf_filter_coeff451_b,rf_filter_coeff452_a, rf_filter_coeff452_b,
    rf_filter_coeff453_a, rf_filter_coeff453_b,rf_filter_coeff454_a, rf_filter_coeff454_b,rf_filter_coeff455_a, rf_filter_coeff455_b,rf_filter_coeff456_a, rf_filter_coeff456_b,
    rf_filter_coeff457_a, rf_filter_coeff457_b,rf_filter_coeff458_a, rf_filter_coeff458_b,rf_filter_coeff459_a, rf_filter_coeff459_b,rf_filter_coeff460_a, rf_filter_coeff460_b,
    rf_filter_coeff461_a, rf_filter_coeff461_b,rf_filter_coeff462_a, rf_filter_coeff462_b,rf_filter_coeff463_a, rf_filter_coeff463_b,rf_filter_coeff464_a, rf_filter_coeff464_b,
    rf_filter_coeff465_a, rf_filter_coeff465_b,rf_filter_coeff466_a, rf_filter_coeff466_b,rf_filter_coeff467_a, rf_filter_coeff467_b,rf_filter_coeff468_a, rf_filter_coeff468_b,
    rf_filter_coeff469_a, rf_filter_coeff469_b,rf_filter_coeff470_a, rf_filter_coeff470_b,rf_filter_coeff471_a, rf_filter_coeff471_b,rf_filter_coeff472_a, rf_filter_coeff472_b,
    rf_filter_coeff473_a, rf_filter_coeff473_b,rf_filter_coeff474_a, rf_filter_coeff474_b,rf_filter_coeff475_a, rf_filter_coeff475_b,rf_filter_coeff476_a, rf_filter_coeff476_b,
    rf_filter_coeff477_a, rf_filter_coeff477_b,rf_filter_coeff478_a, rf_filter_coeff478_b,rf_filter_coeff479_a, rf_filter_coeff479_b,rf_filter_coeff480_a, rf_filter_coeff480_b,
    rf_filter_coeff481_a, rf_filter_coeff481_b,rf_filter_coeff482_a, rf_filter_coeff482_b,rf_filter_coeff483_a, rf_filter_coeff483_b,rf_filter_coeff484_a, rf_filter_coeff484_b,
    rf_filter_coeff485_a, rf_filter_coeff485_b,rf_filter_coeff486_a, rf_filter_coeff486_b,rf_filter_coeff487_a, rf_filter_coeff487_b,rf_filter_coeff488_a, rf_filter_coeff488_b,
    rf_filter_coeff489_a, rf_filter_coeff489_b,rf_filter_coeff490_a, rf_filter_coeff490_b,rf_filter_coeff491_a, rf_filter_coeff491_b,rf_filter_coeff492_a, rf_filter_coeff492_b,
    rf_filter_coeff493_a, rf_filter_coeff493_b,rf_filter_coeff494_a, rf_filter_coeff494_b,rf_filter_coeff495_a, rf_filter_coeff495_b,rf_filter_coeff496_a, rf_filter_coeff496_b,
    rf_filter_coeff497_a, rf_filter_coeff497_b,rf_filter_coeff498_a, rf_filter_coeff498_b,rf_filter_coeff499_a, rf_filter_coeff499_b,rf_filter_coeff500_a, rf_filter_coeff500_b,
    rf_filter_coeff501_a, rf_filter_coeff501_b,rf_filter_coeff502_a, rf_filter_coeff502_b,rf_filter_coeff503_a, rf_filter_coeff503_b,rf_filter_coeff504_a, rf_filter_coeff504_b,
    rf_filter_coeff505_a, rf_filter_coeff505_b,rf_filter_coeff506_a, rf_filter_coeff506_b,rf_filter_coeff507_a, rf_filter_coeff507_b,rf_filter_coeff508_a, rf_filter_coeff508_b,
    rf_filter_coeff509_a, rf_filter_coeff509_b,rf_filter_coeff510_a, rf_filter_coeff510_b,rf_filter_coeff511_a, rf_filter_coeff511_b;
    
    input										clk;
    input										rden;
    input		    [8:0]					    rdptr;
    output	        [15:0]                      rddata;

    localparam	                                DEPTH = 511;        //2^9 = 512
    localparam	                                WIDTH = 15; 

    wire	        [WIDTH:0]                   ram [DEPTH:0];
    reg	            [WIDTH:0]                   rddata;	


    assign ram[0] = {rf_filter_coeff0_b, rf_filter_coeff0_a};
    assign ram[1] = {rf_filter_coeff1_b, rf_filter_coeff1_a};
    assign ram[2] = {rf_filter_coeff2_b, rf_filter_coeff2_a};
    assign ram[3] = {rf_filter_coeff3_b, rf_filter_coeff3_a};
    assign ram[4] = {rf_filter_coeff4_b, rf_filter_coeff4_a};
    assign ram[5] = {rf_filter_coeff5_b, rf_filter_coeff5_a};
    assign ram[6] = {rf_filter_coeff6_b, rf_filter_coeff6_a};
    assign ram[7] = {rf_filter_coeff7_b, rf_filter_coeff7_a};
    assign ram[8] = {rf_filter_coeff8_b, rf_filter_coeff8_a};
    assign ram[9] = {rf_filter_coeff9_b, rf_filter_coeff9_a};
    assign ram[10] = {rf_filter_coeff10_b, rf_filter_coeff10_a};
    assign ram[11] = {rf_filter_coeff11_b, rf_filter_coeff11_a};
    assign ram[12] = {rf_filter_coeff12_b, rf_filter_coeff12_a};
    assign ram[13] = {rf_filter_coeff13_b, rf_filter_coeff13_a};
    assign ram[14] = {rf_filter_coeff14_b, rf_filter_coeff14_a};
    assign ram[15] = {rf_filter_coeff15_b, rf_filter_coeff15_a};
    assign ram[16] = {rf_filter_coeff16_b, rf_filter_coeff16_a};
    assign ram[17] = {rf_filter_coeff17_b, rf_filter_coeff17_a};
    assign ram[18] = {rf_filter_coeff18_b, rf_filter_coeff18_a};
    assign ram[19] = {rf_filter_coeff19_b, rf_filter_coeff19_a};
    assign ram[20] = {rf_filter_coeff20_b, rf_filter_coeff20_a};
    assign ram[21] = {rf_filter_coeff21_b, rf_filter_coeff21_a};
    assign ram[22] = {rf_filter_coeff22_b, rf_filter_coeff22_a};
    assign ram[23] = {rf_filter_coeff23_b, rf_filter_coeff23_a};
    assign ram[24] = {rf_filter_coeff24_b, rf_filter_coeff24_a};
    assign ram[25] = {rf_filter_coeff25_b, rf_filter_coeff25_a};
    assign ram[26] = {rf_filter_coeff26_b, rf_filter_coeff26_a};
    assign ram[27] = {rf_filter_coeff27_b, rf_filter_coeff27_a};
    assign ram[28] = {rf_filter_coeff28_b, rf_filter_coeff28_a};
    assign ram[29] = {rf_filter_coeff29_b, rf_filter_coeff29_a};
    assign ram[30] = {rf_filter_coeff30_b, rf_filter_coeff30_a};
    assign ram[31] = {rf_filter_coeff31_b, rf_filter_coeff31_a};
    assign ram[32] = {rf_filter_coeff32_b, rf_filter_coeff32_a};
    assign ram[33] = {rf_filter_coeff33_b, rf_filter_coeff33_a};
    assign ram[34] = {rf_filter_coeff34_b, rf_filter_coeff34_a};
    assign ram[35] = {rf_filter_coeff35_b, rf_filter_coeff35_a};
    assign ram[36] = {rf_filter_coeff36_b, rf_filter_coeff36_a};
    assign ram[37] = {rf_filter_coeff37_b, rf_filter_coeff37_a};
    assign ram[38] = {rf_filter_coeff38_b, rf_filter_coeff38_a};
    assign ram[39] = {rf_filter_coeff39_b, rf_filter_coeff39_a};
    assign ram[40] = {rf_filter_coeff40_b, rf_filter_coeff40_a};
    assign ram[41] = {rf_filter_coeff41_b, rf_filter_coeff41_a};
    assign ram[42] = {rf_filter_coeff42_b, rf_filter_coeff42_a};
    assign ram[43] = {rf_filter_coeff43_b, rf_filter_coeff43_a};
    assign ram[44] = {rf_filter_coeff44_b, rf_filter_coeff44_a};
    assign ram[45] = {rf_filter_coeff45_b, rf_filter_coeff45_a};
    assign ram[46] = {rf_filter_coeff46_b, rf_filter_coeff46_a};
    assign ram[47] = {rf_filter_coeff47_b, rf_filter_coeff47_a};
    assign ram[48] = {rf_filter_coeff48_b, rf_filter_coeff48_a};
    assign ram[49] = {rf_filter_coeff49_b, rf_filter_coeff49_a};
    assign ram[50] = {rf_filter_coeff50_b, rf_filter_coeff50_a};
    assign ram[51] = {rf_filter_coeff51_b, rf_filter_coeff51_a};
    assign ram[52] = {rf_filter_coeff52_b, rf_filter_coeff52_a};
    assign ram[53] = {rf_filter_coeff53_b, rf_filter_coeff53_a};
    assign ram[54] = {rf_filter_coeff54_b, rf_filter_coeff54_a};
    assign ram[55] = {rf_filter_coeff55_b, rf_filter_coeff55_a};
    assign ram[56] = {rf_filter_coeff56_b, rf_filter_coeff56_a};
    assign ram[57] = {rf_filter_coeff57_b, rf_filter_coeff57_a};
    assign ram[58] = {rf_filter_coeff58_b, rf_filter_coeff58_a};
    assign ram[59] = {rf_filter_coeff59_b, rf_filter_coeff59_a};
    assign ram[60] = {rf_filter_coeff60_b, rf_filter_coeff60_a};
    assign ram[61] = {rf_filter_coeff61_b, rf_filter_coeff61_a};
    assign ram[62] = {rf_filter_coeff62_b, rf_filter_coeff62_a};
    assign ram[63] = {rf_filter_coeff63_b, rf_filter_coeff63_a};
    assign ram[64] = {rf_filter_coeff64_b, rf_filter_coeff64_a};
    assign ram[65] = {rf_filter_coeff65_b, rf_filter_coeff65_a};
    assign ram[66] = {rf_filter_coeff66_b, rf_filter_coeff66_a};
    assign ram[67] = {rf_filter_coeff67_b, rf_filter_coeff67_a};
    assign ram[68] = {rf_filter_coeff68_b, rf_filter_coeff68_a};
    assign ram[69] = {rf_filter_coeff69_b, rf_filter_coeff69_a};
    assign ram[70] = {rf_filter_coeff70_b, rf_filter_coeff70_a};
    assign ram[71] = {rf_filter_coeff71_b, rf_filter_coeff71_a};
    assign ram[72] = {rf_filter_coeff72_b, rf_filter_coeff72_a};
    assign ram[73] = {rf_filter_coeff73_b, rf_filter_coeff73_a};
    assign ram[74] = {rf_filter_coeff74_b, rf_filter_coeff74_a};
    assign ram[75] = {rf_filter_coeff75_b, rf_filter_coeff75_a};
    assign ram[76] = {rf_filter_coeff76_b, rf_filter_coeff76_a};
    assign ram[77] = {rf_filter_coeff77_b, rf_filter_coeff77_a};
    assign ram[78] = {rf_filter_coeff78_b, rf_filter_coeff78_a};
    assign ram[79] = {rf_filter_coeff79_b, rf_filter_coeff79_a};
    assign ram[80] = {rf_filter_coeff80_b, rf_filter_coeff80_a};
    assign ram[81] = {rf_filter_coeff81_b, rf_filter_coeff81_a};
    assign ram[82] = {rf_filter_coeff82_b, rf_filter_coeff82_a};
    assign ram[83] = {rf_filter_coeff83_b, rf_filter_coeff83_a};
    assign ram[84] = {rf_filter_coeff84_b, rf_filter_coeff84_a};
    assign ram[85] = {rf_filter_coeff85_b, rf_filter_coeff85_a};
    assign ram[86] = {rf_filter_coeff86_b, rf_filter_coeff86_a};
    assign ram[87] = {rf_filter_coeff87_b, rf_filter_coeff87_a};
    assign ram[88] = {rf_filter_coeff88_b, rf_filter_coeff88_a};
    assign ram[89] = {rf_filter_coeff89_b, rf_filter_coeff89_a};
    assign ram[90] = {rf_filter_coeff90_b, rf_filter_coeff90_a};
    assign ram[91] = {rf_filter_coeff91_b, rf_filter_coeff91_a};
    assign ram[92] = {rf_filter_coeff92_b, rf_filter_coeff92_a};
    assign ram[93] = {rf_filter_coeff93_b, rf_filter_coeff93_a};
    assign ram[94] = {rf_filter_coeff94_b, rf_filter_coeff94_a};
    assign ram[95] = {rf_filter_coeff95_b, rf_filter_coeff95_a};
    assign ram[96] = {rf_filter_coeff96_b, rf_filter_coeff96_a};
    assign ram[97] = {rf_filter_coeff97_b, rf_filter_coeff97_a};
    assign ram[98] = {rf_filter_coeff98_b, rf_filter_coeff98_a};
    assign ram[99] = {rf_filter_coeff99_b, rf_filter_coeff99_a};
    assign ram[100] = {rf_filter_coeff100_b, rf_filter_coeff100_a};
    assign ram[101] = {rf_filter_coeff101_b, rf_filter_coeff101_a};
    assign ram[102] = {rf_filter_coeff102_b, rf_filter_coeff102_a};
    assign ram[103] = {rf_filter_coeff103_b, rf_filter_coeff103_a};
    assign ram[104] = {rf_filter_coeff104_b, rf_filter_coeff104_a};
    assign ram[105] = {rf_filter_coeff105_b, rf_filter_coeff105_a};
    assign ram[106] = {rf_filter_coeff106_b, rf_filter_coeff106_a};
    assign ram[107] = {rf_filter_coeff107_b, rf_filter_coeff107_a};
    assign ram[108] = {rf_filter_coeff108_b, rf_filter_coeff108_a};
    assign ram[109] = {rf_filter_coeff109_b, rf_filter_coeff109_a};
    assign ram[110] = {rf_filter_coeff110_b, rf_filter_coeff110_a};
    assign ram[111] = {rf_filter_coeff111_b, rf_filter_coeff111_a};
    assign ram[112] = {rf_filter_coeff112_b, rf_filter_coeff112_a};
    assign ram[113] = {rf_filter_coeff113_b, rf_filter_coeff113_a};
    assign ram[114] = {rf_filter_coeff114_b, rf_filter_coeff114_a};
    assign ram[115] = {rf_filter_coeff115_b, rf_filter_coeff115_a};
    assign ram[116] = {rf_filter_coeff116_b, rf_filter_coeff116_a};
    assign ram[117] = {rf_filter_coeff117_b, rf_filter_coeff117_a};
    assign ram[118] = {rf_filter_coeff118_b, rf_filter_coeff118_a};
    assign ram[119] = {rf_filter_coeff119_b, rf_filter_coeff119_a};
    assign ram[120] = {rf_filter_coeff120_b, rf_filter_coeff120_a};
    assign ram[121] = {rf_filter_coeff121_b, rf_filter_coeff121_a};
    assign ram[122] = {rf_filter_coeff122_b, rf_filter_coeff122_a};
    assign ram[123] = {rf_filter_coeff123_b, rf_filter_coeff123_a};
    assign ram[124] = {rf_filter_coeff124_b, rf_filter_coeff124_a};
    assign ram[125] = {rf_filter_coeff125_b, rf_filter_coeff125_a};
    assign ram[126] = {rf_filter_coeff126_b, rf_filter_coeff126_a};
    assign ram[127] = {rf_filter_coeff127_b, rf_filter_coeff127_a};
    assign ram[128] = {rf_filter_coeff128_b, rf_filter_coeff128_a};
    assign ram[129] = {rf_filter_coeff129_b, rf_filter_coeff129_a};
    assign ram[130] = {rf_filter_coeff130_b, rf_filter_coeff130_a};
    assign ram[131] = {rf_filter_coeff131_b, rf_filter_coeff131_a};
    assign ram[132] = {rf_filter_coeff132_b, rf_filter_coeff132_a};
    assign ram[133] = {rf_filter_coeff133_b, rf_filter_coeff133_a};
    assign ram[134] = {rf_filter_coeff134_b, rf_filter_coeff134_a};
    assign ram[135] = {rf_filter_coeff135_b, rf_filter_coeff135_a};
    assign ram[136] = {rf_filter_coeff136_b, rf_filter_coeff136_a};
    assign ram[137] = {rf_filter_coeff137_b, rf_filter_coeff137_a};
    assign ram[138] = {rf_filter_coeff138_b, rf_filter_coeff138_a};
    assign ram[139] = {rf_filter_coeff139_b, rf_filter_coeff139_a};
    assign ram[140] = {rf_filter_coeff140_b, rf_filter_coeff140_a};
    assign ram[141] = {rf_filter_coeff141_b, rf_filter_coeff141_a};
    assign ram[142] = {rf_filter_coeff142_b, rf_filter_coeff142_a};
    assign ram[143] = {rf_filter_coeff143_b, rf_filter_coeff143_a};
    assign ram[144] = {rf_filter_coeff144_b, rf_filter_coeff144_a};
    assign ram[145] = {rf_filter_coeff145_b, rf_filter_coeff145_a};
    assign ram[146] = {rf_filter_coeff146_b, rf_filter_coeff146_a};
    assign ram[147] = {rf_filter_coeff147_b, rf_filter_coeff147_a};
    assign ram[148] = {rf_filter_coeff148_b, rf_filter_coeff148_a};
    assign ram[149] = {rf_filter_coeff149_b, rf_filter_coeff149_a};
    assign ram[150] = {rf_filter_coeff150_b, rf_filter_coeff150_a};
    assign ram[151] = {rf_filter_coeff151_b, rf_filter_coeff151_a};
    assign ram[152] = {rf_filter_coeff152_b, rf_filter_coeff152_a};
    assign ram[153] = {rf_filter_coeff153_b, rf_filter_coeff153_a};
    assign ram[154] = {rf_filter_coeff154_b, rf_filter_coeff154_a};
    assign ram[155] = {rf_filter_coeff155_b, rf_filter_coeff155_a};
    assign ram[156] = {rf_filter_coeff156_b, rf_filter_coeff156_a};
    assign ram[157] = {rf_filter_coeff157_b, rf_filter_coeff157_a};
    assign ram[158] = {rf_filter_coeff158_b, rf_filter_coeff158_a};
    assign ram[159] = {rf_filter_coeff159_b, rf_filter_coeff159_a};
    assign ram[160] = {rf_filter_coeff160_b, rf_filter_coeff160_a};
    assign ram[161] = {rf_filter_coeff161_b, rf_filter_coeff161_a};
    assign ram[162] = {rf_filter_coeff162_b, rf_filter_coeff162_a};
    assign ram[163] = {rf_filter_coeff163_b, rf_filter_coeff163_a};
    assign ram[164] = {rf_filter_coeff164_b, rf_filter_coeff164_a};
    assign ram[165] = {rf_filter_coeff165_b, rf_filter_coeff165_a};
    assign ram[166] = {rf_filter_coeff166_b, rf_filter_coeff166_a};
    assign ram[167] = {rf_filter_coeff167_b, rf_filter_coeff167_a};
    assign ram[168] = {rf_filter_coeff168_b, rf_filter_coeff168_a};
    assign ram[169] = {rf_filter_coeff169_b, rf_filter_coeff169_a};
    assign ram[170] = {rf_filter_coeff170_b, rf_filter_coeff170_a};
    assign ram[171] = {rf_filter_coeff171_b, rf_filter_coeff171_a};
    assign ram[172] = {rf_filter_coeff172_b, rf_filter_coeff172_a};
    assign ram[173] = {rf_filter_coeff173_b, rf_filter_coeff173_a};
    assign ram[174] = {rf_filter_coeff174_b, rf_filter_coeff174_a};
    assign ram[175] = {rf_filter_coeff175_b, rf_filter_coeff175_a};
    assign ram[176] = {rf_filter_coeff176_b, rf_filter_coeff176_a};
    assign ram[177] = {rf_filter_coeff177_b, rf_filter_coeff177_a};
    assign ram[178] = {rf_filter_coeff178_b, rf_filter_coeff178_a};
    assign ram[179] = {rf_filter_coeff179_b, rf_filter_coeff179_a};
    assign ram[180] = {rf_filter_coeff180_b, rf_filter_coeff180_a};
    assign ram[181] = {rf_filter_coeff181_b, rf_filter_coeff181_a};
    assign ram[182] = {rf_filter_coeff182_b, rf_filter_coeff182_a};
    assign ram[183] = {rf_filter_coeff183_b, rf_filter_coeff183_a};
    assign ram[184] = {rf_filter_coeff184_b, rf_filter_coeff184_a};
    assign ram[185] = {rf_filter_coeff185_b, rf_filter_coeff185_a};
    assign ram[186] = {rf_filter_coeff186_b, rf_filter_coeff186_a};
    assign ram[187] = {rf_filter_coeff187_b, rf_filter_coeff187_a};
    assign ram[188] = {rf_filter_coeff188_b, rf_filter_coeff188_a};
    assign ram[189] = {rf_filter_coeff189_b, rf_filter_coeff189_a};
    assign ram[190] = {rf_filter_coeff190_b, rf_filter_coeff190_a};
    assign ram[191] = {rf_filter_coeff191_b, rf_filter_coeff191_a};
    assign ram[192] = {rf_filter_coeff192_b, rf_filter_coeff192_a};
    assign ram[193] = {rf_filter_coeff193_b, rf_filter_coeff193_a};
    assign ram[194] = {rf_filter_coeff194_b, rf_filter_coeff194_a};
    assign ram[195] = {rf_filter_coeff195_b, rf_filter_coeff195_a};
    assign ram[196] = {rf_filter_coeff196_b, rf_filter_coeff196_a};
    assign ram[197] = {rf_filter_coeff197_b, rf_filter_coeff197_a};
    assign ram[198] = {rf_filter_coeff198_b, rf_filter_coeff198_a};
    assign ram[199] = {rf_filter_coeff199_b, rf_filter_coeff199_a};
    assign ram[200] = {rf_filter_coeff200_b, rf_filter_coeff200_a};
    assign ram[201] = {rf_filter_coeff201_b, rf_filter_coeff201_a};
    assign ram[202] = {rf_filter_coeff202_b, rf_filter_coeff202_a};
    assign ram[203] = {rf_filter_coeff203_b, rf_filter_coeff203_a};
    assign ram[204] = {rf_filter_coeff204_b, rf_filter_coeff204_a};
    assign ram[205] = {rf_filter_coeff205_b, rf_filter_coeff205_a};
    assign ram[206] = {rf_filter_coeff206_b, rf_filter_coeff206_a};
    assign ram[207] = {rf_filter_coeff207_b, rf_filter_coeff207_a};
    assign ram[208] = {rf_filter_coeff208_b, rf_filter_coeff208_a};
    assign ram[209] = {rf_filter_coeff209_b, rf_filter_coeff209_a};
    assign ram[210] = {rf_filter_coeff210_b, rf_filter_coeff210_a};
    assign ram[211] = {rf_filter_coeff211_b, rf_filter_coeff211_a};
    assign ram[212] = {rf_filter_coeff212_b, rf_filter_coeff212_a};
    assign ram[213] = {rf_filter_coeff213_b, rf_filter_coeff213_a};
    assign ram[214] = {rf_filter_coeff214_b, rf_filter_coeff214_a};
    assign ram[215] = {rf_filter_coeff215_b, rf_filter_coeff215_a};
    assign ram[216] = {rf_filter_coeff216_b, rf_filter_coeff216_a};
    assign ram[217] = {rf_filter_coeff217_b, rf_filter_coeff217_a};
    assign ram[218] = {rf_filter_coeff218_b, rf_filter_coeff218_a};
    assign ram[219] = {rf_filter_coeff219_b, rf_filter_coeff219_a};
    assign ram[220] = {rf_filter_coeff220_b, rf_filter_coeff220_a};
    assign ram[221] = {rf_filter_coeff221_b, rf_filter_coeff221_a};
    assign ram[222] = {rf_filter_coeff222_b, rf_filter_coeff222_a};
    assign ram[223] = {rf_filter_coeff223_b, rf_filter_coeff223_a};
    assign ram[224] = {rf_filter_coeff224_b, rf_filter_coeff224_a};
    assign ram[225] = {rf_filter_coeff225_b, rf_filter_coeff225_a};
    assign ram[226] = {rf_filter_coeff226_b, rf_filter_coeff226_a};
    assign ram[227] = {rf_filter_coeff227_b, rf_filter_coeff227_a};
    assign ram[228] = {rf_filter_coeff228_b, rf_filter_coeff228_a};
    assign ram[229] = {rf_filter_coeff229_b, rf_filter_coeff229_a};
    assign ram[230] = {rf_filter_coeff230_b, rf_filter_coeff230_a};
    assign ram[231] = {rf_filter_coeff231_b, rf_filter_coeff231_a};
    assign ram[232] = {rf_filter_coeff232_b, rf_filter_coeff232_a};
    assign ram[233] = {rf_filter_coeff233_b, rf_filter_coeff233_a};
    assign ram[234] = {rf_filter_coeff234_b, rf_filter_coeff234_a};
    assign ram[235] = {rf_filter_coeff235_b, rf_filter_coeff235_a};
    assign ram[236] = {rf_filter_coeff236_b, rf_filter_coeff236_a};
    assign ram[237] = {rf_filter_coeff237_b, rf_filter_coeff237_a};
    assign ram[238] = {rf_filter_coeff238_b, rf_filter_coeff238_a};
    assign ram[239] = {rf_filter_coeff239_b, rf_filter_coeff239_a};
    assign ram[240] = {rf_filter_coeff240_b, rf_filter_coeff240_a};
    assign ram[241] = {rf_filter_coeff241_b, rf_filter_coeff241_a};
    assign ram[242] = {rf_filter_coeff242_b, rf_filter_coeff242_a};
    assign ram[243] = {rf_filter_coeff243_b, rf_filter_coeff243_a};
    assign ram[244] = {rf_filter_coeff244_b, rf_filter_coeff244_a};
    assign ram[245] = {rf_filter_coeff245_b, rf_filter_coeff245_a};
    assign ram[246] = {rf_filter_coeff246_b, rf_filter_coeff246_a};
    assign ram[247] = {rf_filter_coeff247_b, rf_filter_coeff247_a};
    assign ram[248] = {rf_filter_coeff248_b, rf_filter_coeff248_a};
    assign ram[249] = {rf_filter_coeff249_b, rf_filter_coeff249_a};
    assign ram[250] = {rf_filter_coeff250_b, rf_filter_coeff250_a};
    assign ram[251] = {rf_filter_coeff251_b, rf_filter_coeff251_a};
    assign ram[252] = {rf_filter_coeff252_b, rf_filter_coeff252_a};
    assign ram[253] = {rf_filter_coeff253_b, rf_filter_coeff253_a};
    assign ram[254] = {rf_filter_coeff254_b, rf_filter_coeff254_a};
    assign ram[255] = {rf_filter_coeff255_b, rf_filter_coeff255_a};
    assign ram[256] = {rf_filter_coeff256_b, rf_filter_coeff256_a};
    assign ram[257] = {rf_filter_coeff257_b, rf_filter_coeff257_a};
    assign ram[258] = {rf_filter_coeff258_b, rf_filter_coeff258_a};
    assign ram[259] = {rf_filter_coeff259_b, rf_filter_coeff259_a};
    assign ram[260] = {rf_filter_coeff260_b, rf_filter_coeff260_a};
    assign ram[261] = {rf_filter_coeff261_b, rf_filter_coeff261_a};
    assign ram[262] = {rf_filter_coeff262_b, rf_filter_coeff262_a};
    assign ram[263] = {rf_filter_coeff263_b, rf_filter_coeff263_a};
    assign ram[264] = {rf_filter_coeff264_b, rf_filter_coeff264_a};
    assign ram[265] = {rf_filter_coeff265_b, rf_filter_coeff265_a};
    assign ram[266] = {rf_filter_coeff266_b, rf_filter_coeff266_a};
    assign ram[267] = {rf_filter_coeff267_b, rf_filter_coeff267_a};
    assign ram[268] = {rf_filter_coeff268_b, rf_filter_coeff268_a};
    assign ram[269] = {rf_filter_coeff269_b, rf_filter_coeff269_a};
    assign ram[270] = {rf_filter_coeff270_b, rf_filter_coeff270_a};
    assign ram[271] = {rf_filter_coeff271_b, rf_filter_coeff271_a};
    assign ram[272] = {rf_filter_coeff272_b, rf_filter_coeff272_a};
    assign ram[273] = {rf_filter_coeff273_b, rf_filter_coeff273_a};
    assign ram[274] = {rf_filter_coeff274_b, rf_filter_coeff274_a};
    assign ram[275] = {rf_filter_coeff275_b, rf_filter_coeff275_a};
    assign ram[276] = {rf_filter_coeff276_b, rf_filter_coeff276_a};
    assign ram[277] = {rf_filter_coeff277_b, rf_filter_coeff277_a};
    assign ram[278] = {rf_filter_coeff278_b, rf_filter_coeff278_a};
    assign ram[279] = {rf_filter_coeff279_b, rf_filter_coeff279_a};
    assign ram[280] = {rf_filter_coeff280_b, rf_filter_coeff280_a};
    assign ram[281] = {rf_filter_coeff281_b, rf_filter_coeff281_a};
    assign ram[282] = {rf_filter_coeff282_b, rf_filter_coeff282_a};
    assign ram[283] = {rf_filter_coeff283_b, rf_filter_coeff283_a};
    assign ram[284] = {rf_filter_coeff284_b, rf_filter_coeff284_a};
    assign ram[285] = {rf_filter_coeff285_b, rf_filter_coeff285_a};
    assign ram[286] = {rf_filter_coeff286_b, rf_filter_coeff286_a};
    assign ram[287] = {rf_filter_coeff287_b, rf_filter_coeff287_a};
    assign ram[288] = {rf_filter_coeff288_b, rf_filter_coeff288_a};
    assign ram[289] = {rf_filter_coeff289_b, rf_filter_coeff289_a};
    assign ram[290] = {rf_filter_coeff290_b, rf_filter_coeff290_a};
    assign ram[291] = {rf_filter_coeff291_b, rf_filter_coeff291_a};
    assign ram[292] = {rf_filter_coeff292_b, rf_filter_coeff292_a};
    assign ram[293] = {rf_filter_coeff293_b, rf_filter_coeff293_a};
    assign ram[294] = {rf_filter_coeff294_b, rf_filter_coeff294_a};
    assign ram[295] = {rf_filter_coeff295_b, rf_filter_coeff295_a};
    assign ram[296] = {rf_filter_coeff296_b, rf_filter_coeff296_a};
    assign ram[297] = {rf_filter_coeff297_b, rf_filter_coeff297_a};
    assign ram[298] = {rf_filter_coeff298_b, rf_filter_coeff298_a};
    assign ram[299] = {rf_filter_coeff299_b, rf_filter_coeff299_a};
    assign ram[300] = {rf_filter_coeff300_b, rf_filter_coeff300_a};
    assign ram[301] = {rf_filter_coeff301_b, rf_filter_coeff301_a};
    assign ram[302] = {rf_filter_coeff302_b, rf_filter_coeff302_a};
    assign ram[303] = {rf_filter_coeff303_b, rf_filter_coeff303_a};
    assign ram[304] = {rf_filter_coeff304_b, rf_filter_coeff304_a};
    assign ram[305] = {rf_filter_coeff305_b, rf_filter_coeff305_a};
    assign ram[306] = {rf_filter_coeff306_b, rf_filter_coeff306_a};
    assign ram[307] = {rf_filter_coeff307_b, rf_filter_coeff307_a};
    assign ram[308] = {rf_filter_coeff308_b, rf_filter_coeff308_a};
    assign ram[309] = {rf_filter_coeff309_b, rf_filter_coeff309_a};
    assign ram[310] = {rf_filter_coeff310_b, rf_filter_coeff310_a};
    assign ram[311] = {rf_filter_coeff311_b, rf_filter_coeff311_a};
    assign ram[312] = {rf_filter_coeff312_b, rf_filter_coeff312_a};
    assign ram[313] = {rf_filter_coeff313_b, rf_filter_coeff313_a};
    assign ram[314] = {rf_filter_coeff314_b, rf_filter_coeff314_a};
    assign ram[315] = {rf_filter_coeff315_b, rf_filter_coeff315_a};
    assign ram[316] = {rf_filter_coeff316_b, rf_filter_coeff316_a};
    assign ram[317] = {rf_filter_coeff317_b, rf_filter_coeff317_a};
    assign ram[318] = {rf_filter_coeff318_b, rf_filter_coeff318_a};
    assign ram[319] = {rf_filter_coeff319_b, rf_filter_coeff319_a};
    assign ram[320] = {rf_filter_coeff320_b, rf_filter_coeff320_a};
    assign ram[321] = {rf_filter_coeff321_b, rf_filter_coeff321_a};
    assign ram[322] = {rf_filter_coeff322_b, rf_filter_coeff322_a};
    assign ram[323] = {rf_filter_coeff323_b, rf_filter_coeff323_a};
    assign ram[324] = {rf_filter_coeff324_b, rf_filter_coeff324_a};
    assign ram[325] = {rf_filter_coeff325_b, rf_filter_coeff325_a};
    assign ram[326] = {rf_filter_coeff326_b, rf_filter_coeff326_a};
    assign ram[327] = {rf_filter_coeff327_b, rf_filter_coeff327_a};
    assign ram[328] = {rf_filter_coeff328_b, rf_filter_coeff328_a};
    assign ram[329] = {rf_filter_coeff329_b, rf_filter_coeff329_a};
    assign ram[330] = {rf_filter_coeff330_b, rf_filter_coeff330_a};
    assign ram[331] = {rf_filter_coeff331_b, rf_filter_coeff331_a};
    assign ram[332] = {rf_filter_coeff332_b, rf_filter_coeff332_a};
    assign ram[333] = {rf_filter_coeff333_b, rf_filter_coeff333_a};
    assign ram[334] = {rf_filter_coeff334_b, rf_filter_coeff334_a};
    assign ram[335] = {rf_filter_coeff335_b, rf_filter_coeff335_a};
    assign ram[336] = {rf_filter_coeff336_b, rf_filter_coeff336_a};
    assign ram[337] = {rf_filter_coeff337_b, rf_filter_coeff337_a};
    assign ram[338] = {rf_filter_coeff338_b, rf_filter_coeff338_a};
    assign ram[339] = {rf_filter_coeff339_b, rf_filter_coeff339_a};
    assign ram[340] = {rf_filter_coeff340_b, rf_filter_coeff340_a};
    assign ram[341] = {rf_filter_coeff341_b, rf_filter_coeff341_a};
    assign ram[342] = {rf_filter_coeff342_b, rf_filter_coeff342_a};
    assign ram[343] = {rf_filter_coeff343_b, rf_filter_coeff343_a};
    assign ram[344] = {rf_filter_coeff344_b, rf_filter_coeff344_a};
    assign ram[345] = {rf_filter_coeff345_b, rf_filter_coeff345_a};
    assign ram[346] = {rf_filter_coeff346_b, rf_filter_coeff346_a};
    assign ram[347] = {rf_filter_coeff347_b, rf_filter_coeff347_a};
    assign ram[348] = {rf_filter_coeff348_b, rf_filter_coeff348_a};
    assign ram[349] = {rf_filter_coeff349_b, rf_filter_coeff349_a};
    assign ram[350] = {rf_filter_coeff350_b, rf_filter_coeff350_a};
    assign ram[351] = {rf_filter_coeff351_b, rf_filter_coeff351_a};
    assign ram[352] = {rf_filter_coeff352_b, rf_filter_coeff352_a};
    assign ram[353] = {rf_filter_coeff353_b, rf_filter_coeff353_a};
    assign ram[354] = {rf_filter_coeff354_b, rf_filter_coeff354_a};
    assign ram[355] = {rf_filter_coeff355_b, rf_filter_coeff355_a};
    assign ram[356] = {rf_filter_coeff356_b, rf_filter_coeff356_a};
    assign ram[357] = {rf_filter_coeff357_b, rf_filter_coeff357_a};
    assign ram[358] = {rf_filter_coeff358_b, rf_filter_coeff358_a};
    assign ram[359] = {rf_filter_coeff359_b, rf_filter_coeff359_a};
    assign ram[360] = {rf_filter_coeff360_b, rf_filter_coeff360_a};
    assign ram[361] = {rf_filter_coeff361_b, rf_filter_coeff361_a};
    assign ram[362] = {rf_filter_coeff362_b, rf_filter_coeff362_a};
    assign ram[363] = {rf_filter_coeff363_b, rf_filter_coeff363_a};
    assign ram[364] = {rf_filter_coeff364_b, rf_filter_coeff364_a};
    assign ram[365] = {rf_filter_coeff365_b, rf_filter_coeff365_a};
    assign ram[366] = {rf_filter_coeff366_b, rf_filter_coeff366_a};
    assign ram[367] = {rf_filter_coeff367_b, rf_filter_coeff367_a};
    assign ram[368] = {rf_filter_coeff368_b, rf_filter_coeff368_a};
    assign ram[369] = {rf_filter_coeff369_b, rf_filter_coeff369_a};
    assign ram[370] = {rf_filter_coeff370_b, rf_filter_coeff370_a};
    assign ram[371] = {rf_filter_coeff371_b, rf_filter_coeff371_a};
    assign ram[372] = {rf_filter_coeff372_b, rf_filter_coeff372_a};
    assign ram[373] = {rf_filter_coeff373_b, rf_filter_coeff373_a};
    assign ram[374] = {rf_filter_coeff374_b, rf_filter_coeff374_a};
    assign ram[375] = {rf_filter_coeff375_b, rf_filter_coeff375_a};
    assign ram[376] = {rf_filter_coeff376_b, rf_filter_coeff376_a};
    assign ram[377] = {rf_filter_coeff377_b, rf_filter_coeff377_a};
    assign ram[378] = {rf_filter_coeff378_b, rf_filter_coeff378_a};
    assign ram[379] = {rf_filter_coeff379_b, rf_filter_coeff379_a};
    assign ram[380] = {rf_filter_coeff380_b, rf_filter_coeff380_a};
    assign ram[381] = {rf_filter_coeff381_b, rf_filter_coeff381_a};
    assign ram[382] = {rf_filter_coeff382_b, rf_filter_coeff382_a};
    assign ram[383] = {rf_filter_coeff383_b, rf_filter_coeff383_a};
    assign ram[384] = {rf_filter_coeff384_b, rf_filter_coeff384_a};
    assign ram[385] = {rf_filter_coeff385_b, rf_filter_coeff385_a};
    assign ram[386] = {rf_filter_coeff386_b, rf_filter_coeff386_a};
    assign ram[387] = {rf_filter_coeff387_b, rf_filter_coeff387_a};
    assign ram[388] = {rf_filter_coeff388_b, rf_filter_coeff388_a};
    assign ram[389] = {rf_filter_coeff389_b, rf_filter_coeff389_a};
    assign ram[390] = {rf_filter_coeff390_b, rf_filter_coeff390_a};
    assign ram[391] = {rf_filter_coeff391_b, rf_filter_coeff391_a};
    assign ram[392] = {rf_filter_coeff392_b, rf_filter_coeff392_a};
    assign ram[393] = {rf_filter_coeff393_b, rf_filter_coeff393_a};
    assign ram[394] = {rf_filter_coeff394_b, rf_filter_coeff394_a};
    assign ram[395] = {rf_filter_coeff395_b, rf_filter_coeff395_a};
    assign ram[396] = {rf_filter_coeff396_b, rf_filter_coeff396_a};
    assign ram[397] = {rf_filter_coeff397_b, rf_filter_coeff397_a};
    assign ram[398] = {rf_filter_coeff398_b, rf_filter_coeff398_a};
    assign ram[399] = {rf_filter_coeff399_b, rf_filter_coeff399_a};
    assign ram[400] = {rf_filter_coeff400_b, rf_filter_coeff400_a};
    assign ram[401] = {rf_filter_coeff401_b, rf_filter_coeff401_a};
    assign ram[402] = {rf_filter_coeff402_b, rf_filter_coeff402_a};
    assign ram[403] = {rf_filter_coeff403_b, rf_filter_coeff403_a};
    assign ram[404] = {rf_filter_coeff404_b, rf_filter_coeff404_a};
    assign ram[405] = {rf_filter_coeff405_b, rf_filter_coeff405_a};
    assign ram[406] = {rf_filter_coeff406_b, rf_filter_coeff406_a};
    assign ram[407] = {rf_filter_coeff407_b, rf_filter_coeff407_a};
    assign ram[408] = {rf_filter_coeff408_b, rf_filter_coeff408_a};
    assign ram[409] = {rf_filter_coeff409_b, rf_filter_coeff409_a};
    assign ram[410] = {rf_filter_coeff410_b, rf_filter_coeff410_a};
    assign ram[411] = {rf_filter_coeff411_b, rf_filter_coeff411_a};
    assign ram[412] = {rf_filter_coeff412_b, rf_filter_coeff412_a};
    assign ram[413] = {rf_filter_coeff413_b, rf_filter_coeff413_a};
    assign ram[414] = {rf_filter_coeff414_b, rf_filter_coeff414_a};
    assign ram[415] = {rf_filter_coeff415_b, rf_filter_coeff415_a};
    assign ram[416] = {rf_filter_coeff416_b, rf_filter_coeff416_a};
    assign ram[417] = {rf_filter_coeff417_b, rf_filter_coeff417_a};
    assign ram[418] = {rf_filter_coeff418_b, rf_filter_coeff418_a};
    assign ram[419] = {rf_filter_coeff419_b, rf_filter_coeff419_a};
    assign ram[420] = {rf_filter_coeff420_b, rf_filter_coeff420_a};
    assign ram[421] = {rf_filter_coeff421_b, rf_filter_coeff421_a};
    assign ram[422] = {rf_filter_coeff422_b, rf_filter_coeff422_a};
    assign ram[423] = {rf_filter_coeff423_b, rf_filter_coeff423_a};
    assign ram[424] = {rf_filter_coeff424_b, rf_filter_coeff424_a};
    assign ram[425] = {rf_filter_coeff425_b, rf_filter_coeff425_a};
    assign ram[426] = {rf_filter_coeff426_b, rf_filter_coeff426_a};
    assign ram[427] = {rf_filter_coeff427_b, rf_filter_coeff427_a};
    assign ram[428] = {rf_filter_coeff428_b, rf_filter_coeff428_a};
    assign ram[429] = {rf_filter_coeff429_b, rf_filter_coeff429_a};
    assign ram[430] = {rf_filter_coeff430_b, rf_filter_coeff430_a};
    assign ram[431] = {rf_filter_coeff431_b, rf_filter_coeff431_a};
    assign ram[432] = {rf_filter_coeff432_b, rf_filter_coeff432_a};
    assign ram[433] = {rf_filter_coeff433_b, rf_filter_coeff433_a};
    assign ram[434] = {rf_filter_coeff434_b, rf_filter_coeff434_a};
    assign ram[435] = {rf_filter_coeff435_b, rf_filter_coeff435_a};
    assign ram[436] = {rf_filter_coeff436_b, rf_filter_coeff436_a};
    assign ram[437] = {rf_filter_coeff437_b, rf_filter_coeff437_a};
    assign ram[438] = {rf_filter_coeff438_b, rf_filter_coeff438_a};
    assign ram[439] = {rf_filter_coeff439_b, rf_filter_coeff439_a};
    assign ram[440] = {rf_filter_coeff440_b, rf_filter_coeff440_a};
    assign ram[441] = {rf_filter_coeff441_b, rf_filter_coeff441_a};
    assign ram[442] = {rf_filter_coeff442_b, rf_filter_coeff442_a};
    assign ram[443] = {rf_filter_coeff443_b, rf_filter_coeff443_a};
    assign ram[444] = {rf_filter_coeff444_b, rf_filter_coeff444_a};
    assign ram[445] = {rf_filter_coeff445_b, rf_filter_coeff445_a};
    assign ram[446] = {rf_filter_coeff446_b, rf_filter_coeff446_a};
    assign ram[447] = {rf_filter_coeff447_b, rf_filter_coeff447_a};
    assign ram[448] = {rf_filter_coeff448_b, rf_filter_coeff448_a};
    assign ram[449] = {rf_filter_coeff449_b, rf_filter_coeff449_a};
    assign ram[450] = {rf_filter_coeff450_b, rf_filter_coeff450_a};
    assign ram[451] = {rf_filter_coeff451_b, rf_filter_coeff451_a};
    assign ram[452] = {rf_filter_coeff452_b, rf_filter_coeff452_a};
    assign ram[453] = {rf_filter_coeff453_b, rf_filter_coeff453_a};
    assign ram[454] = {rf_filter_coeff454_b, rf_filter_coeff454_a};
    assign ram[455] = {rf_filter_coeff455_b, rf_filter_coeff455_a};
    assign ram[456] = {rf_filter_coeff456_b, rf_filter_coeff456_a};
    assign ram[457] = {rf_filter_coeff457_b, rf_filter_coeff457_a};
    assign ram[458] = {rf_filter_coeff458_b, rf_filter_coeff458_a};
    assign ram[459] = {rf_filter_coeff459_b, rf_filter_coeff459_a};
    assign ram[460] = {rf_filter_coeff460_b, rf_filter_coeff460_a};
    assign ram[461] = {rf_filter_coeff461_b, rf_filter_coeff461_a};
    assign ram[462] = {rf_filter_coeff462_b, rf_filter_coeff462_a};
    assign ram[463] = {rf_filter_coeff463_b, rf_filter_coeff463_a};
    assign ram[464] = {rf_filter_coeff464_b, rf_filter_coeff464_a};
    assign ram[465] = {rf_filter_coeff465_b, rf_filter_coeff465_a};
    assign ram[466] = {rf_filter_coeff466_b, rf_filter_coeff466_a};
    assign ram[467] = {rf_filter_coeff467_b, rf_filter_coeff467_a};
    assign ram[468] = {rf_filter_coeff468_b, rf_filter_coeff468_a};
    assign ram[469] = {rf_filter_coeff469_b, rf_filter_coeff469_a};
    assign ram[470] = {rf_filter_coeff470_b, rf_filter_coeff470_a};
    assign ram[471] = {rf_filter_coeff471_b, rf_filter_coeff471_a};
    assign ram[472] = {rf_filter_coeff472_b, rf_filter_coeff472_a};
    assign ram[473] = {rf_filter_coeff473_b, rf_filter_coeff473_a};
    assign ram[474] = {rf_filter_coeff474_b, rf_filter_coeff474_a};
    assign ram[475] = {rf_filter_coeff475_b, rf_filter_coeff475_a};
    assign ram[476] = {rf_filter_coeff476_b, rf_filter_coeff476_a};
    assign ram[477] = {rf_filter_coeff477_b, rf_filter_coeff477_a};
    assign ram[478] = {rf_filter_coeff478_b, rf_filter_coeff478_a};
    assign ram[479] = {rf_filter_coeff479_b, rf_filter_coeff479_a};
    assign ram[480] = {rf_filter_coeff480_b, rf_filter_coeff480_a};
    assign ram[481] = {rf_filter_coeff481_b, rf_filter_coeff481_a};
    assign ram[482] = {rf_filter_coeff482_b, rf_filter_coeff482_a};
    assign ram[483] = {rf_filter_coeff483_b, rf_filter_coeff483_a};
    assign ram[484] = {rf_filter_coeff484_b, rf_filter_coeff484_a};
    assign ram[485] = {rf_filter_coeff485_b, rf_filter_coeff485_a};
    assign ram[486] = {rf_filter_coeff486_b, rf_filter_coeff486_a};
    assign ram[487] = {rf_filter_coeff487_b, rf_filter_coeff487_a};
    assign ram[488] = {rf_filter_coeff488_b, rf_filter_coeff488_a};
    assign ram[489] = {rf_filter_coeff489_b, rf_filter_coeff489_a};
    assign ram[490] = {rf_filter_coeff490_b, rf_filter_coeff490_a};
    assign ram[491] = {rf_filter_coeff491_b, rf_filter_coeff491_a};
    assign ram[492] = {rf_filter_coeff492_b, rf_filter_coeff492_a};
    assign ram[493] = {rf_filter_coeff493_b, rf_filter_coeff493_a};
    assign ram[494] = {rf_filter_coeff494_b, rf_filter_coeff494_a};
    assign ram[495] = {rf_filter_coeff495_b, rf_filter_coeff495_a};
    assign ram[496] = {rf_filter_coeff496_b, rf_filter_coeff496_a};
    assign ram[497] = {rf_filter_coeff497_b, rf_filter_coeff497_a};
    assign ram[498] = {rf_filter_coeff498_b, rf_filter_coeff498_a};
    assign ram[499] = {rf_filter_coeff499_b, rf_filter_coeff499_a};
    assign ram[500] = {rf_filter_coeff500_b, rf_filter_coeff500_a};
    assign ram[501] = {rf_filter_coeff501_b, rf_filter_coeff501_a};
    assign ram[502] = {rf_filter_coeff502_b, rf_filter_coeff502_a};
    assign ram[503] = {rf_filter_coeff503_b, rf_filter_coeff503_a};
    assign ram[504] = {rf_filter_coeff504_b, rf_filter_coeff504_a};
    assign ram[505] = {rf_filter_coeff505_b, rf_filter_coeff505_a};
    assign ram[506] = {rf_filter_coeff506_b, rf_filter_coeff506_a};
    assign ram[507] = {rf_filter_coeff507_b, rf_filter_coeff507_a};
    assign ram[508] = {rf_filter_coeff508_b, rf_filter_coeff508_a};
    assign ram[509] = {rf_filter_coeff509_b, rf_filter_coeff509_a};
    assign ram[510] = {rf_filter_coeff510_b, rf_filter_coeff510_a};
    assign ram[511] = {rf_filter_coeff511_b, rf_filter_coeff511_a};


    always @(posedge clk)
    begin
        if(rden)
            rddata <= ram[rdptr];
    end
    
endmodule
