`timescale 1ns / 1ps

module filter(clk, rstb, aud_in, aud_in_rts, aud_in_rtr, aud_out, aud_out_rts,aud_out_rtr, rf_filter_shift, rf_filter_clip_en, trig_filter_ovf_flag_clear, ro_filter_ovf_flag,
rf_filter_coeff0_a, rf_filter_coeff0_b,rf_filter_coeff1_a, rf_filter_coeff1_b,rf_filter_coeff2_a, rf_filter_coeff2_b,rf_filter_coeff3_a, rf_filter_coeff3_b,rf_filter_coeff4_a, rf_filter_coeff4_b,rf_filter_coeff5_a, rf_filter_coeff5_b,rf_filter_coeff6_a, rf_filter_coeff6_b,rf_filter_coeff7_a, rf_filter_coeff7_b,rf_filter_coeff8_a, rf_filter_coeff8_b,rf_filter_coeff9_a, rf_filter_coeff9_b,rf_filter_coeff10_a, rf_filter_coeff10_b,rf_filter_coeff11_a, rf_filter_coeff11_b,rf_filter_coeff12_a, rf_filter_coeff12_b,rf_filter_coeff13_a, rf_filter_coeff13_b,rf_filter_coeff14_a, rf_filter_coeff14_b,rf_filter_coeff15_a, rf_filter_coeff15_b,rf_filter_coeff16_a, rf_filter_coeff16_b,rf_filter_coeff17_a, rf_filter_coeff17_b,rf_filter_coeff18_a, rf_filter_coeff18_b,rf_filter_coeff19_a, rf_filter_coeff19_b,rf_filter_coeff20_a, rf_filter_coeff20_b,rf_filter_coeff21_a, rf_filter_coeff21_b,rf_filter_coeff22_a, rf_filter_coeff22_b,rf_filter_coeff23_a, rf_filter_coeff23_b,rf_filter_coeff24_a, rf_filter_coeff24_b,rf_filter_coeff25_a, rf_filter_coeff25_b,rf_filter_coeff26_a, rf_filter_coeff26_b,rf_filter_coeff27_a, rf_filter_coeff27_b,rf_filter_coeff28_a, rf_filter_coeff28_b,rf_filter_coeff29_a, rf_filter_coeff29_b,rf_filter_coeff30_a, rf_filter_coeff30_b,rf_filter_coeff31_a, rf_filter_coeff31_b,rf_filter_coeff32_a, rf_filter_coeff32_b,rf_filter_coeff33_a, rf_filter_coeff33_b,rf_filter_coeff34_a, rf_filter_coeff34_b,rf_filter_coeff35_a, rf_filter_coeff35_b,rf_filter_coeff36_a, rf_filter_coeff36_b,rf_filter_coeff37_a, rf_filter_coeff37_b,rf_filter_coeff38_a, rf_filter_coeff38_b,rf_filter_coeff39_a, rf_filter_coeff39_b,rf_filter_coeff40_a, rf_filter_coeff40_b,rf_filter_coeff41_a, rf_filter_coeff41_b,rf_filter_coeff42_a, rf_filter_coeff42_b,rf_filter_coeff43_a, rf_filter_coeff43_b,rf_filter_coeff44_a, rf_filter_coeff44_b,rf_filter_coeff45_a, rf_filter_coeff45_b,rf_filter_coeff46_a, rf_filter_coeff46_b,rf_filter_coeff47_a, rf_filter_coeff47_b,rf_filter_coeff48_a, rf_filter_coeff48_b,rf_filter_coeff49_a, rf_filter_coeff49_b,rf_filter_coeff50_a, rf_filter_coeff50_b,rf_filter_coeff51_a, rf_filter_coeff51_b,rf_filter_coeff52_a, rf_filter_coeff52_b,rf_filter_coeff53_a, rf_filter_coeff53_b,rf_filter_coeff54_a, rf_filter_coeff54_b,rf_filter_coeff55_a, rf_filter_coeff55_b,rf_filter_coeff56_a, rf_filter_coeff56_b,rf_filter_coeff57_a, rf_filter_coeff57_b,rf_filter_coeff58_a, rf_filter_coeff58_b,rf_filter_coeff59_a, rf_filter_coeff59_b,rf_filter_coeff60_a, rf_filter_coeff60_b,rf_filter_coeff61_a, rf_filter_coeff61_b,rf_filter_coeff62_a, rf_filter_coeff62_b,rf_filter_coeff63_a, rf_filter_coeff63_b,rf_filter_coeff64_a, rf_filter_coeff64_b,rf_filter_coeff65_a, rf_filter_coeff65_b,rf_filter_coeff66_a, rf_filter_coeff66_b,rf_filter_coeff67_a, rf_filter_coeff67_b,rf_filter_coeff68_a, rf_filter_coeff68_b,rf_filter_coeff69_a, rf_filter_coeff69_b,rf_filter_coeff70_a, rf_filter_coeff70_b,rf_filter_coeff71_a, rf_filter_coeff71_b,rf_filter_coeff72_a, rf_filter_coeff72_b,rf_filter_coeff73_a, rf_filter_coeff73_b,rf_filter_coeff74_a, rf_filter_coeff74_b,rf_filter_coeff75_a, rf_filter_coeff75_b,rf_filter_coeff76_a, rf_filter_coeff76_b,rf_filter_coeff77_a, rf_filter_coeff77_b,rf_filter_coeff78_a, rf_filter_coeff78_b,rf_filter_coeff79_a, rf_filter_coeff79_b,rf_filter_coeff80_a, rf_filter_coeff80_b,rf_filter_coeff81_a, rf_filter_coeff81_b,rf_filter_coeff82_a, rf_filter_coeff82_b,rf_filter_coeff83_a, rf_filter_coeff83_b,rf_filter_coeff84_a, rf_filter_coeff84_b,rf_filter_coeff85_a, rf_filter_coeff85_b,rf_filter_coeff86_a, rf_filter_coeff86_b,rf_filter_coeff87_a, rf_filter_coeff87_b,rf_filter_coeff88_a, rf_filter_coeff88_b,rf_filter_coeff89_a, rf_filter_coeff89_b,rf_filter_coeff90_a, rf_filter_coeff90_b,rf_filter_coeff91_a, rf_filter_coeff91_b,rf_filter_coeff92_a, rf_filter_coeff92_b,rf_filter_coeff93_a, rf_filter_coeff93_b,rf_filter_coeff94_a, rf_filter_coeff94_b,rf_filter_coeff95_a, rf_filter_coeff95_b,rf_filter_coeff96_a, rf_filter_coeff96_b,rf_filter_coeff97_a, rf_filter_coeff97_b,rf_filter_coeff98_a, rf_filter_coeff98_b,rf_filter_coeff99_a, rf_filter_coeff99_b,rf_filter_coeff100_a, rf_filter_coeff100_b,rf_filter_coeff101_a, rf_filter_coeff101_b,rf_filter_coeff102_a, rf_filter_coeff102_b,rf_filter_coeff103_a, rf_filter_coeff103_b,rf_filter_coeff104_a, rf_filter_coeff104_b,rf_filter_coeff105_a, rf_filter_coeff105_b,rf_filter_coeff106_a, rf_filter_coeff106_b,rf_filter_coeff107_a, rf_filter_coeff107_b,rf_filter_coeff108_a, rf_filter_coeff108_b,rf_filter_coeff109_a, rf_filter_coeff109_b,rf_filter_coeff110_a, rf_filter_coeff110_b,rf_filter_coeff111_a, rf_filter_coeff111_b,rf_filter_coeff112_a, rf_filter_coeff112_b,rf_filter_coeff113_a, rf_filter_coeff113_b,rf_filter_coeff114_a, rf_filter_coeff114_b,rf_filter_coeff115_a, rf_filter_coeff115_b,rf_filter_coeff116_a, rf_filter_coeff116_b,rf_filter_coeff117_a, rf_filter_coeff117_b,rf_filter_coeff118_a, rf_filter_coeff118_b,rf_filter_coeff119_a, rf_filter_coeff119_b,rf_filter_coeff120_a, rf_filter_coeff120_b,rf_filter_coeff121_a, rf_filter_coeff121_b,rf_filter_coeff122_a, rf_filter_coeff122_b,rf_filter_coeff123_a, rf_filter_coeff123_b,rf_filter_coeff124_a, rf_filter_coeff124_b,rf_filter_coeff125_a, rf_filter_coeff125_b,rf_filter_coeff126_a, rf_filter_coeff126_b,rf_filter_coeff127_a, rf_filter_coeff127_b,rf_filter_coeff128_a, rf_filter_coeff128_b,rf_filter_coeff129_a, rf_filter_coeff129_b,rf_filter_coeff130_a, rf_filter_coeff130_b,rf_filter_coeff131_a, rf_filter_coeff131_b,rf_filter_coeff132_a, rf_filter_coeff132_b,rf_filter_coeff133_a, rf_filter_coeff133_b,rf_filter_coeff134_a, rf_filter_coeff134_b,rf_filter_coeff135_a, rf_filter_coeff135_b,rf_filter_coeff136_a, rf_filter_coeff136_b,rf_filter_coeff137_a, rf_filter_coeff137_b,rf_filter_coeff138_a, rf_filter_coeff138_b,rf_filter_coeff139_a, rf_filter_coeff139_b,rf_filter_coeff140_a, rf_filter_coeff140_b,rf_filter_coeff141_a, rf_filter_coeff141_b,rf_filter_coeff142_a, rf_filter_coeff142_b,rf_filter_coeff143_a, rf_filter_coeff143_b,rf_filter_coeff144_a, rf_filter_coeff144_b,rf_filter_coeff145_a, rf_filter_coeff145_b,rf_filter_coeff146_a, rf_filter_coeff146_b,rf_filter_coeff147_a, rf_filter_coeff147_b,rf_filter_coeff148_a, rf_filter_coeff148_b,rf_filter_coeff149_a, rf_filter_coeff149_b,rf_filter_coeff150_a, rf_filter_coeff150_b,rf_filter_coeff151_a, rf_filter_coeff151_b,rf_filter_coeff152_a, rf_filter_coeff152_b,rf_filter_coeff153_a, rf_filter_coeff153_b,rf_filter_coeff154_a, rf_filter_coeff154_b,rf_filter_coeff155_a, rf_filter_coeff155_b,rf_filter_coeff156_a, rf_filter_coeff156_b,rf_filter_coeff157_a, rf_filter_coeff157_b,rf_filter_coeff158_a, rf_filter_coeff158_b,rf_filter_coeff159_a, rf_filter_coeff159_b,rf_filter_coeff160_a, rf_filter_coeff160_b,rf_filter_coeff161_a, rf_filter_coeff161_b,rf_filter_coeff162_a, rf_filter_coeff162_b,rf_filter_coeff163_a, rf_filter_coeff163_b,rf_filter_coeff164_a, rf_filter_coeff164_b,rf_filter_coeff165_a, rf_filter_coeff165_b,rf_filter_coeff166_a, rf_filter_coeff166_b,rf_filter_coeff167_a, rf_filter_coeff167_b,rf_filter_coeff168_a, rf_filter_coeff168_b,rf_filter_coeff169_a, rf_filter_coeff169_b,rf_filter_coeff170_a, rf_filter_coeff170_b,rf_filter_coeff171_a, rf_filter_coeff171_b,rf_filter_coeff172_a, rf_filter_coeff172_b,rf_filter_coeff173_a, rf_filter_coeff173_b,rf_filter_coeff174_a, rf_filter_coeff174_b,rf_filter_coeff175_a, rf_filter_coeff175_b,rf_filter_coeff176_a, rf_filter_coeff176_b,rf_filter_coeff177_a, rf_filter_coeff177_b,rf_filter_coeff178_a, rf_filter_coeff178_b,rf_filter_coeff179_a, rf_filter_coeff179_b,rf_filter_coeff180_a, rf_filter_coeff180_b,rf_filter_coeff181_a, rf_filter_coeff181_b,rf_filter_coeff182_a, rf_filter_coeff182_b,rf_filter_coeff183_a, rf_filter_coeff183_b,rf_filter_coeff184_a, rf_filter_coeff184_b,rf_filter_coeff185_a, rf_filter_coeff185_b,rf_filter_coeff186_a, rf_filter_coeff186_b,rf_filter_coeff187_a, rf_filter_coeff187_b,rf_filter_coeff188_a, rf_filter_coeff188_b,rf_filter_coeff189_a, rf_filter_coeff189_b,rf_filter_coeff190_a, rf_filter_coeff190_b,rf_filter_coeff191_a, rf_filter_coeff191_b,rf_filter_coeff192_a, rf_filter_coeff192_b,rf_filter_coeff193_a, rf_filter_coeff193_b,rf_filter_coeff194_a, rf_filter_coeff194_b,rf_filter_coeff195_a, rf_filter_coeff195_b,rf_filter_coeff196_a, rf_filter_coeff196_b,rf_filter_coeff197_a, rf_filter_coeff197_b,rf_filter_coeff198_a, rf_filter_coeff198_b,rf_filter_coeff199_a, rf_filter_coeff199_b,rf_filter_coeff200_a, rf_filter_coeff200_b,rf_filter_coeff201_a, rf_filter_coeff201_b,rf_filter_coeff202_a, rf_filter_coeff202_b,rf_filter_coeff203_a, rf_filter_coeff203_b,rf_filter_coeff204_a, rf_filter_coeff204_b,rf_filter_coeff205_a, rf_filter_coeff205_b,rf_filter_coeff206_a, rf_filter_coeff206_b,rf_filter_coeff207_a, rf_filter_coeff207_b,rf_filter_coeff208_a, rf_filter_coeff208_b,rf_filter_coeff209_a, rf_filter_coeff209_b,rf_filter_coeff210_a, rf_filter_coeff210_b,rf_filter_coeff211_a, rf_filter_coeff211_b,rf_filter_coeff212_a, rf_filter_coeff212_b,rf_filter_coeff213_a, rf_filter_coeff213_b,rf_filter_coeff214_a, rf_filter_coeff214_b,rf_filter_coeff215_a, rf_filter_coeff215_b,rf_filter_coeff216_a, rf_filter_coeff216_b,rf_filter_coeff217_a, rf_filter_coeff217_b,rf_filter_coeff218_a, rf_filter_coeff218_b,rf_filter_coeff219_a, rf_filter_coeff219_b,rf_filter_coeff220_a, rf_filter_coeff220_b,rf_filter_coeff221_a, rf_filter_coeff221_b,rf_filter_coeff222_a, rf_filter_coeff222_b,rf_filter_coeff223_a, rf_filter_coeff223_b,rf_filter_coeff224_a, rf_filter_coeff224_b,rf_filter_coeff225_a, rf_filter_coeff225_b,rf_filter_coeff226_a, rf_filter_coeff226_b,rf_filter_coeff227_a, rf_filter_coeff227_b,rf_filter_coeff228_a, rf_filter_coeff228_b,rf_filter_coeff229_a, rf_filter_coeff229_b,rf_filter_coeff230_a, rf_filter_coeff230_b,rf_filter_coeff231_a, rf_filter_coeff231_b,rf_filter_coeff232_a, rf_filter_coeff232_b,rf_filter_coeff233_a, rf_filter_coeff233_b,rf_filter_coeff234_a, rf_filter_coeff234_b,rf_filter_coeff235_a, rf_filter_coeff235_b,rf_filter_coeff236_a, rf_filter_coeff236_b,rf_filter_coeff237_a, rf_filter_coeff237_b,rf_filter_coeff238_a, rf_filter_coeff238_b,rf_filter_coeff239_a, rf_filter_coeff239_b,rf_filter_coeff240_a, rf_filter_coeff240_b,rf_filter_coeff241_a, rf_filter_coeff241_b,rf_filter_coeff242_a, rf_filter_coeff242_b,rf_filter_coeff243_a, rf_filter_coeff243_b,rf_filter_coeff244_a, rf_filter_coeff244_b,rf_filter_coeff245_a, rf_filter_coeff245_b,rf_filter_coeff246_a, rf_filter_coeff246_b,rf_filter_coeff247_a, rf_filter_coeff247_b,rf_filter_coeff248_a, rf_filter_coeff248_b,rf_filter_coeff249_a, rf_filter_coeff249_b,rf_filter_coeff250_a, rf_filter_coeff250_b,rf_filter_coeff251_a, rf_filter_coeff251_b,rf_filter_coeff252_a, rf_filter_coeff252_b,rf_filter_coeff253_a, rf_filter_coeff253_b,rf_filter_coeff254_a, rf_filter_coeff254_b,rf_filter_coeff255_a, rf_filter_coeff255_b,rf_filter_coeff256_a, rf_filter_coeff256_b,rf_filter_coeff257_a, rf_filter_coeff257_b,rf_filter_coeff258_a, rf_filter_coeff258_b,rf_filter_coeff259_a, rf_filter_coeff259_b,rf_filter_coeff260_a, rf_filter_coeff260_b,rf_filter_coeff261_a, rf_filter_coeff261_b,rf_filter_coeff262_a, rf_filter_coeff262_b,rf_filter_coeff263_a, rf_filter_coeff263_b,rf_filter_coeff264_a, rf_filter_coeff264_b,rf_filter_coeff265_a, rf_filter_coeff265_b,rf_filter_coeff266_a, rf_filter_coeff266_b,rf_filter_coeff267_a, rf_filter_coeff267_b,rf_filter_coeff268_a, rf_filter_coeff268_b,rf_filter_coeff269_a, rf_filter_coeff269_b,rf_filter_coeff270_a, rf_filter_coeff270_b,rf_filter_coeff271_a, rf_filter_coeff271_b,rf_filter_coeff272_a, rf_filter_coeff272_b,rf_filter_coeff273_a, rf_filter_coeff273_b,rf_filter_coeff274_a, rf_filter_coeff274_b,rf_filter_coeff275_a, rf_filter_coeff275_b,rf_filter_coeff276_a, rf_filter_coeff276_b,rf_filter_coeff277_a, rf_filter_coeff277_b,rf_filter_coeff278_a, rf_filter_coeff278_b,rf_filter_coeff279_a, rf_filter_coeff279_b,rf_filter_coeff280_a, rf_filter_coeff280_b,rf_filter_coeff281_a, rf_filter_coeff281_b,rf_filter_coeff282_a, rf_filter_coeff282_b,rf_filter_coeff283_a, rf_filter_coeff283_b,rf_filter_coeff284_a, rf_filter_coeff284_b,rf_filter_coeff285_a, rf_filter_coeff285_b,rf_filter_coeff286_a, rf_filter_coeff286_b,rf_filter_coeff287_a, rf_filter_coeff287_b,rf_filter_coeff288_a, rf_filter_coeff288_b,rf_filter_coeff289_a, rf_filter_coeff289_b,rf_filter_coeff290_a, rf_filter_coeff290_b,rf_filter_coeff291_a, rf_filter_coeff291_b,rf_filter_coeff292_a, rf_filter_coeff292_b,rf_filter_coeff293_a, rf_filter_coeff293_b,rf_filter_coeff294_a, rf_filter_coeff294_b,rf_filter_coeff295_a, rf_filter_coeff295_b,rf_filter_coeff296_a, rf_filter_coeff296_b,rf_filter_coeff297_a, rf_filter_coeff297_b,rf_filter_coeff298_a, rf_filter_coeff298_b,rf_filter_coeff299_a, rf_filter_coeff299_b,rf_filter_coeff300_a, rf_filter_coeff300_b,rf_filter_coeff301_a, rf_filter_coeff301_b,rf_filter_coeff302_a, rf_filter_coeff302_b,rf_filter_coeff303_a, rf_filter_coeff303_b,rf_filter_coeff304_a, rf_filter_coeff304_b,rf_filter_coeff305_a, rf_filter_coeff305_b,rf_filter_coeff306_a, rf_filter_coeff306_b,rf_filter_coeff307_a, rf_filter_coeff307_b,rf_filter_coeff308_a, rf_filter_coeff308_b,rf_filter_coeff309_a, rf_filter_coeff309_b,rf_filter_coeff310_a, rf_filter_coeff310_b,rf_filter_coeff311_a, rf_filter_coeff311_b,rf_filter_coeff312_a, rf_filter_coeff312_b,rf_filter_coeff313_a, rf_filter_coeff313_b,rf_filter_coeff314_a, rf_filter_coeff314_b,rf_filter_coeff315_a, rf_filter_coeff315_b,rf_filter_coeff316_a, rf_filter_coeff316_b,rf_filter_coeff317_a, rf_filter_coeff317_b,rf_filter_coeff318_a, rf_filter_coeff318_b,rf_filter_coeff319_a, rf_filter_coeff319_b,rf_filter_coeff320_a, rf_filter_coeff320_b,rf_filter_coeff321_a, rf_filter_coeff321_b,rf_filter_coeff322_a, rf_filter_coeff322_b,rf_filter_coeff323_a, rf_filter_coeff323_b,rf_filter_coeff324_a, rf_filter_coeff324_b,rf_filter_coeff325_a, rf_filter_coeff325_b,rf_filter_coeff326_a, rf_filter_coeff326_b,rf_filter_coeff327_a, rf_filter_coeff327_b,rf_filter_coeff328_a, rf_filter_coeff328_b,rf_filter_coeff329_a, rf_filter_coeff329_b,rf_filter_coeff330_a, rf_filter_coeff330_b,rf_filter_coeff331_a, rf_filter_coeff331_b,rf_filter_coeff332_a, rf_filter_coeff332_b,rf_filter_coeff333_a, rf_filter_coeff333_b,rf_filter_coeff334_a, rf_filter_coeff334_b,rf_filter_coeff335_a, rf_filter_coeff335_b,rf_filter_coeff336_a, rf_filter_coeff336_b,rf_filter_coeff337_a, rf_filter_coeff337_b,rf_filter_coeff338_a, rf_filter_coeff338_b,rf_filter_coeff339_a, rf_filter_coeff339_b,rf_filter_coeff340_a, rf_filter_coeff340_b,rf_filter_coeff341_a, rf_filter_coeff341_b,rf_filter_coeff342_a, rf_filter_coeff342_b,rf_filter_coeff343_a, rf_filter_coeff343_b,rf_filter_coeff344_a, rf_filter_coeff344_b,rf_filter_coeff345_a, rf_filter_coeff345_b,rf_filter_coeff346_a, rf_filter_coeff346_b,rf_filter_coeff347_a, rf_filter_coeff347_b,rf_filter_coeff348_a, rf_filter_coeff348_b,rf_filter_coeff349_a, rf_filter_coeff349_b,rf_filter_coeff350_a, rf_filter_coeff350_b,rf_filter_coeff351_a, rf_filter_coeff351_b,rf_filter_coeff352_a, rf_filter_coeff352_b,rf_filter_coeff353_a, rf_filter_coeff353_b,rf_filter_coeff354_a, rf_filter_coeff354_b,rf_filter_coeff355_a, rf_filter_coeff355_b,rf_filter_coeff356_a, rf_filter_coeff356_b,rf_filter_coeff357_a, rf_filter_coeff357_b,rf_filter_coeff358_a, rf_filter_coeff358_b,rf_filter_coeff359_a, rf_filter_coeff359_b,rf_filter_coeff360_a, rf_filter_coeff360_b,rf_filter_coeff361_a, rf_filter_coeff361_b,rf_filter_coeff362_a, rf_filter_coeff362_b,rf_filter_coeff363_a, rf_filter_coeff363_b,rf_filter_coeff364_a, rf_filter_coeff364_b,rf_filter_coeff365_a, rf_filter_coeff365_b,rf_filter_coeff366_a, rf_filter_coeff366_b,rf_filter_coeff367_a, rf_filter_coeff367_b,rf_filter_coeff368_a, rf_filter_coeff368_b,rf_filter_coeff369_a, rf_filter_coeff369_b,rf_filter_coeff370_a, rf_filter_coeff370_b,rf_filter_coeff371_a, rf_filter_coeff371_b,rf_filter_coeff372_a, rf_filter_coeff372_b,rf_filter_coeff373_a, rf_filter_coeff373_b,rf_filter_coeff374_a, rf_filter_coeff374_b,rf_filter_coeff375_a, rf_filter_coeff375_b,rf_filter_coeff376_a, rf_filter_coeff376_b,rf_filter_coeff377_a, rf_filter_coeff377_b,rf_filter_coeff378_a, rf_filter_coeff378_b,rf_filter_coeff379_a, rf_filter_coeff379_b,rf_filter_coeff380_a, rf_filter_coeff380_b,rf_filter_coeff381_a, rf_filter_coeff381_b,rf_filter_coeff382_a, rf_filter_coeff382_b,rf_filter_coeff383_a, rf_filter_coeff383_b,rf_filter_coeff384_a, rf_filter_coeff384_b,rf_filter_coeff385_a, rf_filter_coeff385_b,rf_filter_coeff386_a, rf_filter_coeff386_b,rf_filter_coeff387_a, rf_filter_coeff387_b,rf_filter_coeff388_a, rf_filter_coeff388_b,rf_filter_coeff389_a, rf_filter_coeff389_b,rf_filter_coeff390_a, rf_filter_coeff390_b,rf_filter_coeff391_a, rf_filter_coeff391_b,rf_filter_coeff392_a, rf_filter_coeff392_b,rf_filter_coeff393_a, rf_filter_coeff393_b,rf_filter_coeff394_a, rf_filter_coeff394_b,rf_filter_coeff395_a, rf_filter_coeff395_b,rf_filter_coeff396_a, rf_filter_coeff396_b,rf_filter_coeff397_a, rf_filter_coeff397_b,rf_filter_coeff398_a, rf_filter_coeff398_b,rf_filter_coeff399_a, rf_filter_coeff399_b,rf_filter_coeff400_a, rf_filter_coeff400_b,rf_filter_coeff401_a, rf_filter_coeff401_b,rf_filter_coeff402_a, rf_filter_coeff402_b,rf_filter_coeff403_a, rf_filter_coeff403_b,rf_filter_coeff404_a, rf_filter_coeff404_b,rf_filter_coeff405_a, rf_filter_coeff405_b,rf_filter_coeff406_a, rf_filter_coeff406_b,rf_filter_coeff407_a, rf_filter_coeff407_b,rf_filter_coeff408_a, rf_filter_coeff408_b,rf_filter_coeff409_a, rf_filter_coeff409_b,rf_filter_coeff410_a, rf_filter_coeff410_b,rf_filter_coeff411_a, rf_filter_coeff411_b,rf_filter_coeff412_a, rf_filter_coeff412_b,rf_filter_coeff413_a, rf_filter_coeff413_b,rf_filter_coeff414_a, rf_filter_coeff414_b,rf_filter_coeff415_a, rf_filter_coeff415_b,rf_filter_coeff416_a, rf_filter_coeff416_b,rf_filter_coeff417_a, rf_filter_coeff417_b,rf_filter_coeff418_a, rf_filter_coeff418_b,rf_filter_coeff419_a, rf_filter_coeff419_b,rf_filter_coeff420_a, rf_filter_coeff420_b,rf_filter_coeff421_a, rf_filter_coeff421_b,rf_filter_coeff422_a, rf_filter_coeff422_b,rf_filter_coeff423_a, rf_filter_coeff423_b,rf_filter_coeff424_a, rf_filter_coeff424_b,rf_filter_coeff425_a, rf_filter_coeff425_b,rf_filter_coeff426_a, rf_filter_coeff426_b,rf_filter_coeff427_a, rf_filter_coeff427_b,rf_filter_coeff428_a, rf_filter_coeff428_b,rf_filter_coeff429_a, rf_filter_coeff429_b,rf_filter_coeff430_a, rf_filter_coeff430_b,rf_filter_coeff431_a, rf_filter_coeff431_b,rf_filter_coeff432_a, rf_filter_coeff432_b,rf_filter_coeff433_a, rf_filter_coeff433_b,rf_filter_coeff434_a, rf_filter_coeff434_b,rf_filter_coeff435_a, rf_filter_coeff435_b,rf_filter_coeff436_a, rf_filter_coeff436_b,rf_filter_coeff437_a, rf_filter_coeff437_b,rf_filter_coeff438_a, rf_filter_coeff438_b,rf_filter_coeff439_a, rf_filter_coeff439_b,rf_filter_coeff440_a, rf_filter_coeff440_b,rf_filter_coeff441_a, rf_filter_coeff441_b,rf_filter_coeff442_a, rf_filter_coeff442_b,rf_filter_coeff443_a, rf_filter_coeff443_b,rf_filter_coeff444_a, rf_filter_coeff444_b,rf_filter_coeff445_a, rf_filter_coeff445_b,rf_filter_coeff446_a, rf_filter_coeff446_b,rf_filter_coeff447_a, rf_filter_coeff447_b,rf_filter_coeff448_a, rf_filter_coeff448_b,rf_filter_coeff449_a, rf_filter_coeff449_b,rf_filter_coeff450_a, rf_filter_coeff450_b,rf_filter_coeff451_a, rf_filter_coeff451_b,rf_filter_coeff452_a, rf_filter_coeff452_b,rf_filter_coeff453_a, rf_filter_coeff453_b,rf_filter_coeff454_a, rf_filter_coeff454_b,rf_filter_coeff455_a, rf_filter_coeff455_b,rf_filter_coeff456_a, rf_filter_coeff456_b,rf_filter_coeff457_a, rf_filter_coeff457_b,rf_filter_coeff458_a, rf_filter_coeff458_b,rf_filter_coeff459_a, rf_filter_coeff459_b,rf_filter_coeff460_a, rf_filter_coeff460_b,rf_filter_coeff461_a, rf_filter_coeff461_b,rf_filter_coeff462_a, rf_filter_coeff462_b,rf_filter_coeff463_a, rf_filter_coeff463_b,rf_filter_coeff464_a, rf_filter_coeff464_b,rf_filter_coeff465_a, rf_filter_coeff465_b,rf_filter_coeff466_a, rf_filter_coeff466_b,rf_filter_coeff467_a, rf_filter_coeff467_b,rf_filter_coeff468_a, rf_filter_coeff468_b,rf_filter_coeff469_a, rf_filter_coeff469_b,rf_filter_coeff470_a, rf_filter_coeff470_b,rf_filter_coeff471_a, rf_filter_coeff471_b,rf_filter_coeff472_a, rf_filter_coeff472_b,rf_filter_coeff473_a, rf_filter_coeff473_b,rf_filter_coeff474_a, rf_filter_coeff474_b,rf_filter_coeff475_a, rf_filter_coeff475_b,rf_filter_coeff476_a, rf_filter_coeff476_b,rf_filter_coeff477_a, rf_filter_coeff477_b,rf_filter_coeff478_a, rf_filter_coeff478_b,rf_filter_coeff479_a, rf_filter_coeff479_b,rf_filter_coeff480_a, rf_filter_coeff480_b,rf_filter_coeff481_a, rf_filter_coeff481_b,rf_filter_coeff482_a, rf_filter_coeff482_b,rf_filter_coeff483_a, rf_filter_coeff483_b,rf_filter_coeff484_a, rf_filter_coeff484_b,rf_filter_coeff485_a, rf_filter_coeff485_b,rf_filter_coeff486_a, rf_filter_coeff486_b,rf_filter_coeff487_a, rf_filter_coeff487_b,rf_filter_coeff488_a, rf_filter_coeff488_b,rf_filter_coeff489_a, rf_filter_coeff489_b,rf_filter_coeff490_a, rf_filter_coeff490_b,rf_filter_coeff491_a, rf_filter_coeff491_b,rf_filter_coeff492_a, rf_filter_coeff492_b,rf_filter_coeff493_a, rf_filter_coeff493_b,rf_filter_coeff494_a, rf_filter_coeff494_b,rf_filter_coeff495_a, rf_filter_coeff495_b,rf_filter_coeff496_a, rf_filter_coeff496_b,rf_filter_coeff497_a, rf_filter_coeff497_b,rf_filter_coeff498_a, rf_filter_coeff498_b,rf_filter_coeff499_a, rf_filter_coeff499_b,rf_filter_coeff500_a, rf_filter_coeff500_b,rf_filter_coeff501_a, rf_filter_coeff501_b,rf_filter_coeff502_a, rf_filter_coeff502_b,rf_filter_coeff503_a, rf_filter_coeff503_b,rf_filter_coeff504_a, rf_filter_coeff504_b,rf_filter_coeff505_a, rf_filter_coeff505_b,rf_filter_coeff506_a, rf_filter_coeff506_b,rf_filter_coeff507_a, rf_filter_coeff507_b,rf_filter_coeff508_a, rf_filter_coeff508_b,rf_filter_coeff509_a, rf_filter_coeff509_b,rf_filter_coeff510_a, rf_filter_coeff510_b,rf_filter_coeff511_a, rf_filter_coeff511_b
     );

input 	clk;
input 	rstb;
input 	[31:0] aud_in;
input 	aud_in_rts;
output 	aud_in_rtr;
output 	[31:0] aud_out;
output 	aud_out_rts;
input 	aud_out_rtr;
input 	trig_filter_ovf_flag_clear;
output 	ro_filter_ovf_flag;
input		[2:0] rf_filter_shift;
input		rf_filter_clip_en;
input 	[7:0] rf_filter_coeff0_a, rf_filter_coeff0_b,
rf_filter_coeff1_a, rf_filter_coeff1_b,rf_filter_coeff2_a, rf_filter_coeff2_b,rf_filter_coeff3_a, rf_filter_coeff3_b,rf_filter_coeff4_a, rf_filter_coeff4_b,
rf_filter_coeff5_a, rf_filter_coeff5_b,rf_filter_coeff6_a, rf_filter_coeff6_b,rf_filter_coeff7_a, rf_filter_coeff7_b,rf_filter_coeff8_a, rf_filter_coeff8_b,
rf_filter_coeff9_a, rf_filter_coeff9_b,rf_filter_coeff10_a, rf_filter_coeff10_b,rf_filter_coeff11_a, rf_filter_coeff11_b,rf_filter_coeff12_a, rf_filter_coeff12_b,
rf_filter_coeff13_a, rf_filter_coeff13_b,rf_filter_coeff14_a, rf_filter_coeff14_b,rf_filter_coeff15_a, rf_filter_coeff15_b,rf_filter_coeff16_a, rf_filter_coeff16_b,
rf_filter_coeff17_a, rf_filter_coeff17_b,rf_filter_coeff18_a, rf_filter_coeff18_b,rf_filter_coeff19_a, rf_filter_coeff19_b,rf_filter_coeff20_a, rf_filter_coeff20_b,
rf_filter_coeff21_a, rf_filter_coeff21_b,rf_filter_coeff22_a, rf_filter_coeff22_b,rf_filter_coeff23_a, rf_filter_coeff23_b,rf_filter_coeff24_a, rf_filter_coeff24_b,
rf_filter_coeff25_a, rf_filter_coeff25_b,rf_filter_coeff26_a, rf_filter_coeff26_b,rf_filter_coeff27_a, rf_filter_coeff27_b,rf_filter_coeff28_a, rf_filter_coeff28_b,
rf_filter_coeff29_a, rf_filter_coeff29_b,rf_filter_coeff30_a, rf_filter_coeff30_b,rf_filter_coeff31_a, rf_filter_coeff31_b,rf_filter_coeff32_a, rf_filter_coeff32_b,
rf_filter_coeff33_a, rf_filter_coeff33_b,rf_filter_coeff34_a, rf_filter_coeff34_b,rf_filter_coeff35_a, rf_filter_coeff35_b,rf_filter_coeff36_a, rf_filter_coeff36_b,
rf_filter_coeff37_a, rf_filter_coeff37_b,rf_filter_coeff38_a, rf_filter_coeff38_b,rf_filter_coeff39_a, rf_filter_coeff39_b,rf_filter_coeff40_a, rf_filter_coeff40_b,
rf_filter_coeff41_a, rf_filter_coeff41_b,rf_filter_coeff42_a, rf_filter_coeff42_b,rf_filter_coeff43_a, rf_filter_coeff43_b,rf_filter_coeff44_a, rf_filter_coeff44_b,
rf_filter_coeff45_a, rf_filter_coeff45_b,rf_filter_coeff46_a, rf_filter_coeff46_b,rf_filter_coeff47_a, rf_filter_coeff47_b,rf_filter_coeff48_a, rf_filter_coeff48_b,
rf_filter_coeff49_a, rf_filter_coeff49_b,rf_filter_coeff50_a, rf_filter_coeff50_b,rf_filter_coeff51_a, rf_filter_coeff51_b,rf_filter_coeff52_a, rf_filter_coeff52_b,
rf_filter_coeff53_a, rf_filter_coeff53_b,rf_filter_coeff54_a, rf_filter_coeff54_b,rf_filter_coeff55_a, rf_filter_coeff55_b,rf_filter_coeff56_a, rf_filter_coeff56_b,
rf_filter_coeff57_a, rf_filter_coeff57_b,rf_filter_coeff58_a, rf_filter_coeff58_b,rf_filter_coeff59_a, rf_filter_coeff59_b,rf_filter_coeff60_a, rf_filter_coeff60_b,
rf_filter_coeff61_a, rf_filter_coeff61_b,rf_filter_coeff62_a, rf_filter_coeff62_b,rf_filter_coeff63_a, rf_filter_coeff63_b,rf_filter_coeff64_a, rf_filter_coeff64_b,
rf_filter_coeff65_a, rf_filter_coeff65_b,rf_filter_coeff66_a, rf_filter_coeff66_b,rf_filter_coeff67_a, rf_filter_coeff67_b,rf_filter_coeff68_a, rf_filter_coeff68_b,
rf_filter_coeff69_a, rf_filter_coeff69_b,rf_filter_coeff70_a, rf_filter_coeff70_b,rf_filter_coeff71_a, rf_filter_coeff71_b,rf_filter_coeff72_a, rf_filter_coeff72_b,
rf_filter_coeff73_a, rf_filter_coeff73_b,rf_filter_coeff74_a, rf_filter_coeff74_b,rf_filter_coeff75_a, rf_filter_coeff75_b,rf_filter_coeff76_a, rf_filter_coeff76_b,
rf_filter_coeff77_a, rf_filter_coeff77_b,rf_filter_coeff78_a, rf_filter_coeff78_b,rf_filter_coeff79_a, rf_filter_coeff79_b,rf_filter_coeff80_a, rf_filter_coeff80_b,
rf_filter_coeff81_a, rf_filter_coeff81_b,rf_filter_coeff82_a, rf_filter_coeff82_b,rf_filter_coeff83_a, rf_filter_coeff83_b,rf_filter_coeff84_a, rf_filter_coeff84_b,
rf_filter_coeff85_a, rf_filter_coeff85_b,rf_filter_coeff86_a, rf_filter_coeff86_b,rf_filter_coeff87_a, rf_filter_coeff87_b,rf_filter_coeff88_a, rf_filter_coeff88_b,
rf_filter_coeff89_a, rf_filter_coeff89_b,rf_filter_coeff90_a, rf_filter_coeff90_b,rf_filter_coeff91_a, rf_filter_coeff91_b,rf_filter_coeff92_a, rf_filter_coeff92_b,
rf_filter_coeff93_a, rf_filter_coeff93_b,rf_filter_coeff94_a, rf_filter_coeff94_b,rf_filter_coeff95_a, rf_filter_coeff95_b,rf_filter_coeff96_a, rf_filter_coeff96_b,
rf_filter_coeff97_a, rf_filter_coeff97_b,rf_filter_coeff98_a, rf_filter_coeff98_b,rf_filter_coeff99_a, rf_filter_coeff99_b,rf_filter_coeff100_a, rf_filter_coeff100_b,
rf_filter_coeff101_a, rf_filter_coeff101_b,rf_filter_coeff102_a, rf_filter_coeff102_b,rf_filter_coeff103_a, rf_filter_coeff103_b,rf_filter_coeff104_a, rf_filter_coeff104_b,
rf_filter_coeff105_a, rf_filter_coeff105_b,rf_filter_coeff106_a, rf_filter_coeff106_b,rf_filter_coeff107_a, rf_filter_coeff107_b,rf_filter_coeff108_a, rf_filter_coeff108_b,
rf_filter_coeff109_a, rf_filter_coeff109_b,rf_filter_coeff110_a, rf_filter_coeff110_b,rf_filter_coeff111_a, rf_filter_coeff111_b,rf_filter_coeff112_a, rf_filter_coeff112_b,
rf_filter_coeff113_a, rf_filter_coeff113_b,rf_filter_coeff114_a, rf_filter_coeff114_b,rf_filter_coeff115_a, rf_filter_coeff115_b,rf_filter_coeff116_a, rf_filter_coeff116_b,
rf_filter_coeff117_a, rf_filter_coeff117_b,rf_filter_coeff118_a, rf_filter_coeff118_b,rf_filter_coeff119_a, rf_filter_coeff119_b,rf_filter_coeff120_a, rf_filter_coeff120_b,
rf_filter_coeff121_a, rf_filter_coeff121_b,rf_filter_coeff122_a, rf_filter_coeff122_b,rf_filter_coeff123_a, rf_filter_coeff123_b,rf_filter_coeff124_a, rf_filter_coeff124_b,
rf_filter_coeff125_a, rf_filter_coeff125_b,rf_filter_coeff126_a, rf_filter_coeff126_b,rf_filter_coeff127_a, rf_filter_coeff127_b,rf_filter_coeff128_a, rf_filter_coeff128_b,
rf_filter_coeff129_a, rf_filter_coeff129_b,rf_filter_coeff130_a, rf_filter_coeff130_b,rf_filter_coeff131_a, rf_filter_coeff131_b,rf_filter_coeff132_a, rf_filter_coeff132_b,
rf_filter_coeff133_a, rf_filter_coeff133_b,rf_filter_coeff134_a, rf_filter_coeff134_b,rf_filter_coeff135_a, rf_filter_coeff135_b,rf_filter_coeff136_a, rf_filter_coeff136_b,
rf_filter_coeff137_a, rf_filter_coeff137_b,rf_filter_coeff138_a, rf_filter_coeff138_b,rf_filter_coeff139_a, rf_filter_coeff139_b,rf_filter_coeff140_a, rf_filter_coeff140_b,
rf_filter_coeff141_a, rf_filter_coeff141_b,rf_filter_coeff142_a, rf_filter_coeff142_b,rf_filter_coeff143_a, rf_filter_coeff143_b,rf_filter_coeff144_a, rf_filter_coeff144_b,
rf_filter_coeff145_a, rf_filter_coeff145_b,rf_filter_coeff146_a, rf_filter_coeff146_b,rf_filter_coeff147_a, rf_filter_coeff147_b,rf_filter_coeff148_a, rf_filter_coeff148_b,
rf_filter_coeff149_a, rf_filter_coeff149_b,rf_filter_coeff150_a, rf_filter_coeff150_b,rf_filter_coeff151_a, rf_filter_coeff151_b,rf_filter_coeff152_a, rf_filter_coeff152_b,
rf_filter_coeff153_a, rf_filter_coeff153_b,rf_filter_coeff154_a, rf_filter_coeff154_b,rf_filter_coeff155_a, rf_filter_coeff155_b,rf_filter_coeff156_a, rf_filter_coeff156_b,
rf_filter_coeff157_a, rf_filter_coeff157_b,rf_filter_coeff158_a, rf_filter_coeff158_b,rf_filter_coeff159_a, rf_filter_coeff159_b,rf_filter_coeff160_a, rf_filter_coeff160_b,
rf_filter_coeff161_a, rf_filter_coeff161_b,rf_filter_coeff162_a, rf_filter_coeff162_b,rf_filter_coeff163_a, rf_filter_coeff163_b,rf_filter_coeff164_a, rf_filter_coeff164_b,
rf_filter_coeff165_a, rf_filter_coeff165_b,rf_filter_coeff166_a, rf_filter_coeff166_b,rf_filter_coeff167_a, rf_filter_coeff167_b,rf_filter_coeff168_a, rf_filter_coeff168_b,
rf_filter_coeff169_a, rf_filter_coeff169_b,rf_filter_coeff170_a, rf_filter_coeff170_b,rf_filter_coeff171_a, rf_filter_coeff171_b,rf_filter_coeff172_a, rf_filter_coeff172_b,
rf_filter_coeff173_a, rf_filter_coeff173_b,rf_filter_coeff174_a, rf_filter_coeff174_b,rf_filter_coeff175_a, rf_filter_coeff175_b,rf_filter_coeff176_a, rf_filter_coeff176_b,
rf_filter_coeff177_a, rf_filter_coeff177_b,rf_filter_coeff178_a, rf_filter_coeff178_b,rf_filter_coeff179_a, rf_filter_coeff179_b,rf_filter_coeff180_a, rf_filter_coeff180_b,
rf_filter_coeff181_a, rf_filter_coeff181_b,rf_filter_coeff182_a, rf_filter_coeff182_b,rf_filter_coeff183_a, rf_filter_coeff183_b,rf_filter_coeff184_a, rf_filter_coeff184_b,
rf_filter_coeff185_a, rf_filter_coeff185_b,rf_filter_coeff186_a, rf_filter_coeff186_b,rf_filter_coeff187_a, rf_filter_coeff187_b,rf_filter_coeff188_a, rf_filter_coeff188_b,
rf_filter_coeff189_a, rf_filter_coeff189_b,rf_filter_coeff190_a, rf_filter_coeff190_b,rf_filter_coeff191_a, rf_filter_coeff191_b,rf_filter_coeff192_a, rf_filter_coeff192_b,
rf_filter_coeff193_a, rf_filter_coeff193_b,rf_filter_coeff194_a, rf_filter_coeff194_b,rf_filter_coeff195_a, rf_filter_coeff195_b,rf_filter_coeff196_a, rf_filter_coeff196_b,
rf_filter_coeff197_a, rf_filter_coeff197_b,rf_filter_coeff198_a, rf_filter_coeff198_b,rf_filter_coeff199_a, rf_filter_coeff199_b,rf_filter_coeff200_a, rf_filter_coeff200_b,
rf_filter_coeff201_a, rf_filter_coeff201_b,rf_filter_coeff202_a, rf_filter_coeff202_b,rf_filter_coeff203_a, rf_filter_coeff203_b,rf_filter_coeff204_a, rf_filter_coeff204_b,
rf_filter_coeff205_a, rf_filter_coeff205_b,rf_filter_coeff206_a, rf_filter_coeff206_b,rf_filter_coeff207_a, rf_filter_coeff207_b,rf_filter_coeff208_a, rf_filter_coeff208_b,
rf_filter_coeff209_a, rf_filter_coeff209_b,rf_filter_coeff210_a, rf_filter_coeff210_b,rf_filter_coeff211_a, rf_filter_coeff211_b,rf_filter_coeff212_a, rf_filter_coeff212_b,
rf_filter_coeff213_a, rf_filter_coeff213_b,rf_filter_coeff214_a, rf_filter_coeff214_b,rf_filter_coeff215_a, rf_filter_coeff215_b,rf_filter_coeff216_a, rf_filter_coeff216_b,
rf_filter_coeff217_a, rf_filter_coeff217_b,rf_filter_coeff218_a, rf_filter_coeff218_b,rf_filter_coeff219_a, rf_filter_coeff219_b,rf_filter_coeff220_a, rf_filter_coeff220_b,
rf_filter_coeff221_a, rf_filter_coeff221_b,rf_filter_coeff222_a, rf_filter_coeff222_b,rf_filter_coeff223_a, rf_filter_coeff223_b,rf_filter_coeff224_a, rf_filter_coeff224_b,
rf_filter_coeff225_a, rf_filter_coeff225_b,rf_filter_coeff226_a, rf_filter_coeff226_b,rf_filter_coeff227_a, rf_filter_coeff227_b,rf_filter_coeff228_a, rf_filter_coeff228_b,
rf_filter_coeff229_a, rf_filter_coeff229_b,rf_filter_coeff230_a, rf_filter_coeff230_b,rf_filter_coeff231_a, rf_filter_coeff231_b,rf_filter_coeff232_a, rf_filter_coeff232_b,
rf_filter_coeff233_a, rf_filter_coeff233_b,rf_filter_coeff234_a, rf_filter_coeff234_b,rf_filter_coeff235_a, rf_filter_coeff235_b,rf_filter_coeff236_a, rf_filter_coeff236_b,
rf_filter_coeff237_a, rf_filter_coeff237_b,rf_filter_coeff238_a, rf_filter_coeff238_b,rf_filter_coeff239_a, rf_filter_coeff239_b,rf_filter_coeff240_a, rf_filter_coeff240_b,
rf_filter_coeff241_a, rf_filter_coeff241_b,rf_filter_coeff242_a, rf_filter_coeff242_b,rf_filter_coeff243_a, rf_filter_coeff243_b,rf_filter_coeff244_a, rf_filter_coeff244_b,
rf_filter_coeff245_a, rf_filter_coeff245_b,rf_filter_coeff246_a, rf_filter_coeff246_b,rf_filter_coeff247_a, rf_filter_coeff247_b,rf_filter_coeff248_a, rf_filter_coeff248_b,
rf_filter_coeff249_a, rf_filter_coeff249_b,rf_filter_coeff250_a, rf_filter_coeff250_b,rf_filter_coeff251_a, rf_filter_coeff251_b,rf_filter_coeff252_a, rf_filter_coeff252_b,
rf_filter_coeff253_a, rf_filter_coeff253_b,rf_filter_coeff254_a, rf_filter_coeff254_b,rf_filter_coeff255_a, rf_filter_coeff255_b,rf_filter_coeff256_a, rf_filter_coeff256_b,
rf_filter_coeff257_a, rf_filter_coeff257_b,rf_filter_coeff258_a, rf_filter_coeff258_b,rf_filter_coeff259_a, rf_filter_coeff259_b,rf_filter_coeff260_a, rf_filter_coeff260_b,
rf_filter_coeff261_a, rf_filter_coeff261_b,rf_filter_coeff262_a, rf_filter_coeff262_b,rf_filter_coeff263_a, rf_filter_coeff263_b,rf_filter_coeff264_a, rf_filter_coeff264_b,
rf_filter_coeff265_a, rf_filter_coeff265_b,rf_filter_coeff266_a, rf_filter_coeff266_b,rf_filter_coeff267_a, rf_filter_coeff267_b,rf_filter_coeff268_a, rf_filter_coeff268_b,
rf_filter_coeff269_a, rf_filter_coeff269_b,rf_filter_coeff270_a, rf_filter_coeff270_b,rf_filter_coeff271_a, rf_filter_coeff271_b,rf_filter_coeff272_a, rf_filter_coeff272_b,
rf_filter_coeff273_a, rf_filter_coeff273_b,rf_filter_coeff274_a, rf_filter_coeff274_b,rf_filter_coeff275_a, rf_filter_coeff275_b,rf_filter_coeff276_a, rf_filter_coeff276_b,
rf_filter_coeff277_a, rf_filter_coeff277_b,rf_filter_coeff278_a, rf_filter_coeff278_b,rf_filter_coeff279_a, rf_filter_coeff279_b,rf_filter_coeff280_a, rf_filter_coeff280_b,
rf_filter_coeff281_a, rf_filter_coeff281_b,rf_filter_coeff282_a, rf_filter_coeff282_b,rf_filter_coeff283_a, rf_filter_coeff283_b,rf_filter_coeff284_a, rf_filter_coeff284_b,
rf_filter_coeff285_a, rf_filter_coeff285_b,rf_filter_coeff286_a, rf_filter_coeff286_b,rf_filter_coeff287_a, rf_filter_coeff287_b,rf_filter_coeff288_a, rf_filter_coeff288_b,
rf_filter_coeff289_a, rf_filter_coeff289_b,rf_filter_coeff290_a, rf_filter_coeff290_b,rf_filter_coeff291_a, rf_filter_coeff291_b,rf_filter_coeff292_a, rf_filter_coeff292_b,
rf_filter_coeff293_a, rf_filter_coeff293_b,rf_filter_coeff294_a, rf_filter_coeff294_b,rf_filter_coeff295_a, rf_filter_coeff295_b,rf_filter_coeff296_a, rf_filter_coeff296_b,
rf_filter_coeff297_a, rf_filter_coeff297_b,rf_filter_coeff298_a, rf_filter_coeff298_b,rf_filter_coeff299_a, rf_filter_coeff299_b,rf_filter_coeff300_a, rf_filter_coeff300_b,
rf_filter_coeff301_a, rf_filter_coeff301_b,rf_filter_coeff302_a, rf_filter_coeff302_b,rf_filter_coeff303_a, rf_filter_coeff303_b,rf_filter_coeff304_a, rf_filter_coeff304_b,
rf_filter_coeff305_a, rf_filter_coeff305_b,rf_filter_coeff306_a, rf_filter_coeff306_b,rf_filter_coeff307_a, rf_filter_coeff307_b,rf_filter_coeff308_a, rf_filter_coeff308_b,
rf_filter_coeff309_a, rf_filter_coeff309_b,rf_filter_coeff310_a, rf_filter_coeff310_b,rf_filter_coeff311_a, rf_filter_coeff311_b,rf_filter_coeff312_a, rf_filter_coeff312_b,
rf_filter_coeff313_a, rf_filter_coeff313_b,rf_filter_coeff314_a, rf_filter_coeff314_b,rf_filter_coeff315_a, rf_filter_coeff315_b,rf_filter_coeff316_a, rf_filter_coeff316_b,
rf_filter_coeff317_a, rf_filter_coeff317_b,rf_filter_coeff318_a, rf_filter_coeff318_b,rf_filter_coeff319_a, rf_filter_coeff319_b,rf_filter_coeff320_a, rf_filter_coeff320_b,
rf_filter_coeff321_a, rf_filter_coeff321_b,rf_filter_coeff322_a, rf_filter_coeff322_b,rf_filter_coeff323_a, rf_filter_coeff323_b,rf_filter_coeff324_a, rf_filter_coeff324_b,
rf_filter_coeff325_a, rf_filter_coeff325_b,rf_filter_coeff326_a, rf_filter_coeff326_b,rf_filter_coeff327_a, rf_filter_coeff327_b,rf_filter_coeff328_a, rf_filter_coeff328_b,
rf_filter_coeff329_a, rf_filter_coeff329_b,rf_filter_coeff330_a, rf_filter_coeff330_b,rf_filter_coeff331_a, rf_filter_coeff331_b,rf_filter_coeff332_a, rf_filter_coeff332_b,
rf_filter_coeff333_a, rf_filter_coeff333_b,rf_filter_coeff334_a, rf_filter_coeff334_b,rf_filter_coeff335_a, rf_filter_coeff335_b,rf_filter_coeff336_a, rf_filter_coeff336_b,
rf_filter_coeff337_a, rf_filter_coeff337_b,rf_filter_coeff338_a, rf_filter_coeff338_b,rf_filter_coeff339_a, rf_filter_coeff339_b,rf_filter_coeff340_a, rf_filter_coeff340_b,
rf_filter_coeff341_a, rf_filter_coeff341_b,rf_filter_coeff342_a, rf_filter_coeff342_b,rf_filter_coeff343_a, rf_filter_coeff343_b,rf_filter_coeff344_a, rf_filter_coeff344_b,
rf_filter_coeff345_a, rf_filter_coeff345_b,rf_filter_coeff346_a, rf_filter_coeff346_b,rf_filter_coeff347_a, rf_filter_coeff347_b,rf_filter_coeff348_a, rf_filter_coeff348_b,
rf_filter_coeff349_a, rf_filter_coeff349_b,rf_filter_coeff350_a, rf_filter_coeff350_b,rf_filter_coeff351_a, rf_filter_coeff351_b,rf_filter_coeff352_a, rf_filter_coeff352_b,
rf_filter_coeff353_a, rf_filter_coeff353_b,rf_filter_coeff354_a, rf_filter_coeff354_b,rf_filter_coeff355_a, rf_filter_coeff355_b,rf_filter_coeff356_a, rf_filter_coeff356_b,
rf_filter_coeff357_a, rf_filter_coeff357_b,rf_filter_coeff358_a, rf_filter_coeff358_b,rf_filter_coeff359_a, rf_filter_coeff359_b,rf_filter_coeff360_a, rf_filter_coeff360_b,
rf_filter_coeff361_a, rf_filter_coeff361_b,rf_filter_coeff362_a, rf_filter_coeff362_b,rf_filter_coeff363_a, rf_filter_coeff363_b,rf_filter_coeff364_a, rf_filter_coeff364_b,
rf_filter_coeff365_a, rf_filter_coeff365_b,rf_filter_coeff366_a, rf_filter_coeff366_b,rf_filter_coeff367_a, rf_filter_coeff367_b,rf_filter_coeff368_a, rf_filter_coeff368_b,
rf_filter_coeff369_a, rf_filter_coeff369_b,rf_filter_coeff370_a, rf_filter_coeff370_b,rf_filter_coeff371_a, rf_filter_coeff371_b,rf_filter_coeff372_a, rf_filter_coeff372_b,
rf_filter_coeff373_a, rf_filter_coeff373_b,rf_filter_coeff374_a, rf_filter_coeff374_b,rf_filter_coeff375_a, rf_filter_coeff375_b,rf_filter_coeff376_a, rf_filter_coeff376_b,
rf_filter_coeff377_a, rf_filter_coeff377_b,rf_filter_coeff378_a, rf_filter_coeff378_b,rf_filter_coeff379_a, rf_filter_coeff379_b,rf_filter_coeff380_a, rf_filter_coeff380_b,
rf_filter_coeff381_a, rf_filter_coeff381_b,rf_filter_coeff382_a, rf_filter_coeff382_b,rf_filter_coeff383_a, rf_filter_coeff383_b,rf_filter_coeff384_a, rf_filter_coeff384_b,
rf_filter_coeff385_a, rf_filter_coeff385_b,rf_filter_coeff386_a, rf_filter_coeff386_b,rf_filter_coeff387_a, rf_filter_coeff387_b,rf_filter_coeff388_a, rf_filter_coeff388_b,
rf_filter_coeff389_a, rf_filter_coeff389_b,rf_filter_coeff390_a, rf_filter_coeff390_b,rf_filter_coeff391_a, rf_filter_coeff391_b,rf_filter_coeff392_a, rf_filter_coeff392_b,
rf_filter_coeff393_a, rf_filter_coeff393_b,rf_filter_coeff394_a, rf_filter_coeff394_b,rf_filter_coeff395_a, rf_filter_coeff395_b,rf_filter_coeff396_a, rf_filter_coeff396_b,
rf_filter_coeff397_a, rf_filter_coeff397_b,rf_filter_coeff398_a, rf_filter_coeff398_b,rf_filter_coeff399_a, rf_filter_coeff399_b,rf_filter_coeff400_a, rf_filter_coeff400_b,
rf_filter_coeff401_a, rf_filter_coeff401_b,rf_filter_coeff402_a, rf_filter_coeff402_b,rf_filter_coeff403_a, rf_filter_coeff403_b,rf_filter_coeff404_a, rf_filter_coeff404_b,
rf_filter_coeff405_a, rf_filter_coeff405_b,rf_filter_coeff406_a, rf_filter_coeff406_b,rf_filter_coeff407_a, rf_filter_coeff407_b,rf_filter_coeff408_a, rf_filter_coeff408_b,
rf_filter_coeff409_a, rf_filter_coeff409_b,rf_filter_coeff410_a, rf_filter_coeff410_b,rf_filter_coeff411_a, rf_filter_coeff411_b,rf_filter_coeff412_a, rf_filter_coeff412_b,
rf_filter_coeff413_a, rf_filter_coeff413_b,rf_filter_coeff414_a, rf_filter_coeff414_b,rf_filter_coeff415_a, rf_filter_coeff415_b,rf_filter_coeff416_a, rf_filter_coeff416_b,
rf_filter_coeff417_a, rf_filter_coeff417_b,rf_filter_coeff418_a, rf_filter_coeff418_b,rf_filter_coeff419_a, rf_filter_coeff419_b,rf_filter_coeff420_a, rf_filter_coeff420_b,
rf_filter_coeff421_a, rf_filter_coeff421_b,rf_filter_coeff422_a, rf_filter_coeff422_b,rf_filter_coeff423_a, rf_filter_coeff423_b,rf_filter_coeff424_a, rf_filter_coeff424_b,
rf_filter_coeff425_a, rf_filter_coeff425_b,rf_filter_coeff426_a, rf_filter_coeff426_b,rf_filter_coeff427_a, rf_filter_coeff427_b,rf_filter_coeff428_a, rf_filter_coeff428_b,
rf_filter_coeff429_a, rf_filter_coeff429_b,rf_filter_coeff430_a, rf_filter_coeff430_b,rf_filter_coeff431_a, rf_filter_coeff431_b,rf_filter_coeff432_a, rf_filter_coeff432_b,
rf_filter_coeff433_a, rf_filter_coeff433_b,rf_filter_coeff434_a, rf_filter_coeff434_b,rf_filter_coeff435_a, rf_filter_coeff435_b,rf_filter_coeff436_a, rf_filter_coeff436_b,
rf_filter_coeff437_a, rf_filter_coeff437_b,rf_filter_coeff438_a, rf_filter_coeff438_b,rf_filter_coeff439_a, rf_filter_coeff439_b,rf_filter_coeff440_a, rf_filter_coeff440_b,
rf_filter_coeff441_a, rf_filter_coeff441_b,rf_filter_coeff442_a, rf_filter_coeff442_b,rf_filter_coeff443_a, rf_filter_coeff443_b,rf_filter_coeff444_a, rf_filter_coeff444_b,
rf_filter_coeff445_a, rf_filter_coeff445_b,rf_filter_coeff446_a, rf_filter_coeff446_b,rf_filter_coeff447_a, rf_filter_coeff447_b,rf_filter_coeff448_a, rf_filter_coeff448_b,
rf_filter_coeff449_a, rf_filter_coeff449_b,rf_filter_coeff450_a, rf_filter_coeff450_b,rf_filter_coeff451_a, rf_filter_coeff451_b,rf_filter_coeff452_a, rf_filter_coeff452_b,
rf_filter_coeff453_a, rf_filter_coeff453_b,rf_filter_coeff454_a, rf_filter_coeff454_b,rf_filter_coeff455_a, rf_filter_coeff455_b,rf_filter_coeff456_a, rf_filter_coeff456_b,
rf_filter_coeff457_a, rf_filter_coeff457_b,rf_filter_coeff458_a, rf_filter_coeff458_b,rf_filter_coeff459_a, rf_filter_coeff459_b,rf_filter_coeff460_a, rf_filter_coeff460_b,
rf_filter_coeff461_a, rf_filter_coeff461_b,rf_filter_coeff462_a, rf_filter_coeff462_b,rf_filter_coeff463_a, rf_filter_coeff463_b,rf_filter_coeff464_a, rf_filter_coeff464_b,
rf_filter_coeff465_a, rf_filter_coeff465_b,rf_filter_coeff466_a, rf_filter_coeff466_b,rf_filter_coeff467_a, rf_filter_coeff467_b,rf_filter_coeff468_a, rf_filter_coeff468_b,
rf_filter_coeff469_a, rf_filter_coeff469_b,rf_filter_coeff470_a, rf_filter_coeff470_b,rf_filter_coeff471_a, rf_filter_coeff471_b,rf_filter_coeff472_a, rf_filter_coeff472_b,
rf_filter_coeff473_a, rf_filter_coeff473_b,rf_filter_coeff474_a, rf_filter_coeff474_b,rf_filter_coeff475_a, rf_filter_coeff475_b,rf_filter_coeff476_a, rf_filter_coeff476_b,
rf_filter_coeff477_a, rf_filter_coeff477_b,rf_filter_coeff478_a, rf_filter_coeff478_b,rf_filter_coeff479_a, rf_filter_coeff479_b,rf_filter_coeff480_a, rf_filter_coeff480_b,
rf_filter_coeff481_a, rf_filter_coeff481_b,rf_filter_coeff482_a, rf_filter_coeff482_b,rf_filter_coeff483_a, rf_filter_coeff483_b,rf_filter_coeff484_a, rf_filter_coeff484_b,
rf_filter_coeff485_a, rf_filter_coeff485_b,rf_filter_coeff486_a, rf_filter_coeff486_b,rf_filter_coeff487_a, rf_filter_coeff487_b,rf_filter_coeff488_a, rf_filter_coeff488_b,
rf_filter_coeff489_a, rf_filter_coeff489_b,rf_filter_coeff490_a, rf_filter_coeff490_b,rf_filter_coeff491_a, rf_filter_coeff491_b,rf_filter_coeff492_a, rf_filter_coeff492_b,
rf_filter_coeff493_a, rf_filter_coeff493_b,rf_filter_coeff494_a, rf_filter_coeff494_b,rf_filter_coeff495_a, rf_filter_coeff495_b,rf_filter_coeff496_a, rf_filter_coeff496_b,
rf_filter_coeff497_a, rf_filter_coeff497_b,rf_filter_coeff498_a, rf_filter_coeff498_b,rf_filter_coeff499_a, rf_filter_coeff499_b,rf_filter_coeff500_a, rf_filter_coeff500_b,
rf_filter_coeff501_a, rf_filter_coeff501_b,rf_filter_coeff502_a, rf_filter_coeff502_b,rf_filter_coeff503_a, rf_filter_coeff503_b,rf_filter_coeff504_a, rf_filter_coeff504_b,
rf_filter_coeff505_a, rf_filter_coeff505_b,rf_filter_coeff506_a, rf_filter_coeff506_b,rf_filter_coeff507_a, rf_filter_coeff507_b,rf_filter_coeff508_a, rf_filter_coeff508_b,
rf_filter_coeff509_a, rf_filter_coeff509_b,rf_filter_coeff510_a, rf_filter_coeff510_b,rf_filter_coeff511_a, rf_filter_coeff511_b;

wire 			do_transfer;
wire 			do_multiply_1st;
wire 			do_multiply;
wire[15:0]	rf_filter_coeff;
wire[8:0]	mux_rdptr;			 
wire			mux_re;
wire 			output_signal; 
wire[31:0]	convo_signal;

//assign aud_out = convo_signal[39:8]; 

//***********************************************************************************
filter_stm filter_stm_0 (
    .clk(clk), 
    .rstb(rstb), 
    .filter_aud_in_rts(aud_in_rts), 
    .filter_aud_in_rtr(aud_in_rtr), 
	 .filter_aud_out_rts(aud_out_rts), 
    .filter_aud_out_rtr(aud_out_rtr), 
    .do_transfer(do_transfer), 
    .do_multiply_1st(do_multiply_1st), 
    .do_multiply(do_multiply), 
    .filter_aud_in(aud_in), 
    .filter_aud_out(convo_signal), 
    .rf_filter_coeff(rf_filter_coeff),
	 .rf_shift(rf_filter_shift), 
    .rf_sat(rf_filter_clip_en), 
	 .mux_re(mux_re),
	 .mux_rdptr(mux_rdptr)
    );
	 
	 
	 
//***********************************************************************************

//***********************************************************************************
filter_mux filter_mux_0 (
    .clk(clk), 
    .rden(mux_re), 
    .rdptr(mux_rdptr), 
    .rddata(rf_filter_coeff), 
    .rf_filter_coeff0_a(rf_filter_coeff0_a), 
    .rf_filter_coeff0_b(rf_filter_coeff0_b), 
    .rf_filter_coeff1_a(rf_filter_coeff1_a), 
    .rf_filter_coeff1_b(rf_filter_coeff1_b), 
    .rf_filter_coeff2_a(rf_filter_coeff2_a), 
    .rf_filter_coeff2_b(rf_filter_coeff2_b), 
    .rf_filter_coeff3_a(rf_filter_coeff3_a), 
    .rf_filter_coeff3_b(rf_filter_coeff3_b), 
    .rf_filter_coeff4_a(rf_filter_coeff4_a), 
    .rf_filter_coeff4_b(rf_filter_coeff4_b), 
    .rf_filter_coeff5_a(rf_filter_coeff5_a), 
    .rf_filter_coeff5_b(rf_filter_coeff5_b), 
    .rf_filter_coeff6_a(rf_filter_coeff6_a), 
    .rf_filter_coeff6_b(rf_filter_coeff6_b), 
    .rf_filter_coeff7_a(rf_filter_coeff7_a), 
    .rf_filter_coeff7_b(rf_filter_coeff7_b), 
    .rf_filter_coeff8_a(rf_filter_coeff8_a), 
    .rf_filter_coeff8_b(rf_filter_coeff8_b), 
    .rf_filter_coeff9_a(rf_filter_coeff9_a), 
    .rf_filter_coeff9_b(rf_filter_coeff9_b), 
    .rf_filter_coeff10_a(rf_filter_coeff10_a), 
    .rf_filter_coeff10_b(rf_filter_coeff10_b), 
    .rf_filter_coeff11_a(rf_filter_coeff11_a), 
    .rf_filter_coeff11_b(rf_filter_coeff11_b), 
    .rf_filter_coeff12_a(rf_filter_coeff12_a), 
    .rf_filter_coeff12_b(rf_filter_coeff12_b), 
    .rf_filter_coeff13_a(rf_filter_coeff13_a), 
    .rf_filter_coeff13_b(rf_filter_coeff13_b), 
    .rf_filter_coeff14_a(rf_filter_coeff14_a), 
    .rf_filter_coeff14_b(rf_filter_coeff14_b), 
    .rf_filter_coeff15_a(rf_filter_coeff15_a), 
    .rf_filter_coeff15_b(rf_filter_coeff15_b), 
    .rf_filter_coeff16_a(rf_filter_coeff16_a), 
    .rf_filter_coeff16_b(rf_filter_coeff16_b), 
    .rf_filter_coeff17_a(rf_filter_coeff17_a), 
    .rf_filter_coeff17_b(rf_filter_coeff17_b), 
    .rf_filter_coeff18_a(rf_filter_coeff18_a), 
    .rf_filter_coeff18_b(rf_filter_coeff18_b), 
    .rf_filter_coeff19_a(rf_filter_coeff19_a), 
    .rf_filter_coeff19_b(rf_filter_coeff19_b), 
    .rf_filter_coeff20_a(rf_filter_coeff20_a), 
    .rf_filter_coeff20_b(rf_filter_coeff20_b), 
    .rf_filter_coeff21_a(rf_filter_coeff21_a), 
    .rf_filter_coeff21_b(rf_filter_coeff21_b), 
    .rf_filter_coeff22_a(rf_filter_coeff22_a), 
    .rf_filter_coeff22_b(rf_filter_coeff22_b), 
    .rf_filter_coeff23_a(rf_filter_coeff23_a), 
    .rf_filter_coeff23_b(rf_filter_coeff23_b), 
    .rf_filter_coeff24_a(rf_filter_coeff24_a), 
    .rf_filter_coeff24_b(rf_filter_coeff24_b), 
    .rf_filter_coeff25_a(rf_filter_coeff25_a), 
    .rf_filter_coeff25_b(rf_filter_coeff25_b), 
    .rf_filter_coeff26_a(rf_filter_coeff26_a), 
    .rf_filter_coeff26_b(rf_filter_coeff26_b), 
    .rf_filter_coeff27_a(rf_filter_coeff27_a), 
    .rf_filter_coeff27_b(rf_filter_coeff27_b), 
    .rf_filter_coeff28_a(rf_filter_coeff28_a), 
    .rf_filter_coeff28_b(rf_filter_coeff28_b), 
    .rf_filter_coeff29_a(rf_filter_coeff29_a), 
    .rf_filter_coeff29_b(rf_filter_coeff29_b), 
    .rf_filter_coeff30_a(rf_filter_coeff30_a), 
    .rf_filter_coeff30_b(rf_filter_coeff30_b), 
    .rf_filter_coeff31_a(rf_filter_coeff31_a), 
    .rf_filter_coeff31_b(rf_filter_coeff31_b), 
    .rf_filter_coeff32_a(rf_filter_coeff32_a), 
    .rf_filter_coeff32_b(rf_filter_coeff32_b), 
    .rf_filter_coeff33_a(rf_filter_coeff33_a), 
    .rf_filter_coeff33_b(rf_filter_coeff33_b), 
    .rf_filter_coeff34_a(rf_filter_coeff34_a), 
    .rf_filter_coeff34_b(rf_filter_coeff34_b), 
    .rf_filter_coeff35_a(rf_filter_coeff35_a), 
    .rf_filter_coeff35_b(rf_filter_coeff35_b), 
    .rf_filter_coeff36_a(rf_filter_coeff36_a), 
    .rf_filter_coeff36_b(rf_filter_coeff36_b), 
    .rf_filter_coeff37_a(rf_filter_coeff37_a), 
    .rf_filter_coeff37_b(rf_filter_coeff37_b), 
    .rf_filter_coeff38_a(rf_filter_coeff38_a), 
    .rf_filter_coeff38_b(rf_filter_coeff38_b), 
    .rf_filter_coeff39_a(rf_filter_coeff39_a), 
    .rf_filter_coeff39_b(rf_filter_coeff39_b), 
    .rf_filter_coeff40_a(rf_filter_coeff40_a), 
    .rf_filter_coeff40_b(rf_filter_coeff40_b), 
    .rf_filter_coeff41_a(rf_filter_coeff41_a), 
    .rf_filter_coeff41_b(rf_filter_coeff41_b), 
    .rf_filter_coeff42_a(rf_filter_coeff42_a), 
    .rf_filter_coeff42_b(rf_filter_coeff42_b), 
    .rf_filter_coeff43_a(rf_filter_coeff43_a), 
    .rf_filter_coeff43_b(rf_filter_coeff43_b), 
    .rf_filter_coeff44_a(rf_filter_coeff44_a), 
    .rf_filter_coeff44_b(rf_filter_coeff44_b), 
    .rf_filter_coeff45_a(rf_filter_coeff45_a), 
    .rf_filter_coeff45_b(rf_filter_coeff45_b), 
    .rf_filter_coeff46_a(rf_filter_coeff46_a), 
    .rf_filter_coeff46_b(rf_filter_coeff46_b), 
    .rf_filter_coeff47_a(rf_filter_coeff47_a), 
    .rf_filter_coeff47_b(rf_filter_coeff47_b), 
    .rf_filter_coeff48_a(rf_filter_coeff48_a), 
    .rf_filter_coeff48_b(rf_filter_coeff48_b), 
    .rf_filter_coeff49_a(rf_filter_coeff49_a), 
    .rf_filter_coeff49_b(rf_filter_coeff49_b), 
    .rf_filter_coeff50_a(rf_filter_coeff50_a), 
    .rf_filter_coeff50_b(rf_filter_coeff50_b), 
    .rf_filter_coeff51_a(rf_filter_coeff51_a), 
    .rf_filter_coeff51_b(rf_filter_coeff51_b), 
    .rf_filter_coeff52_a(rf_filter_coeff52_a), 
    .rf_filter_coeff52_b(rf_filter_coeff52_b), 
    .rf_filter_coeff53_a(rf_filter_coeff53_a), 
    .rf_filter_coeff53_b(rf_filter_coeff53_b), 
    .rf_filter_coeff54_a(rf_filter_coeff54_a), 
    .rf_filter_coeff54_b(rf_filter_coeff54_b), 
    .rf_filter_coeff55_a(rf_filter_coeff55_a), 
    .rf_filter_coeff55_b(rf_filter_coeff55_b), 
    .rf_filter_coeff56_a(rf_filter_coeff56_a), 
    .rf_filter_coeff56_b(rf_filter_coeff56_b), 
    .rf_filter_coeff57_a(rf_filter_coeff57_a), 
    .rf_filter_coeff57_b(rf_filter_coeff57_b), 
    .rf_filter_coeff58_a(rf_filter_coeff58_a), 
    .rf_filter_coeff58_b(rf_filter_coeff58_b), 
    .rf_filter_coeff59_a(rf_filter_coeff59_a), 
    .rf_filter_coeff59_b(rf_filter_coeff59_b), 
    .rf_filter_coeff60_a(rf_filter_coeff60_a), 
    .rf_filter_coeff60_b(rf_filter_coeff60_b), 
    .rf_filter_coeff61_a(rf_filter_coeff61_a), 
    .rf_filter_coeff61_b(rf_filter_coeff61_b), 
    .rf_filter_coeff62_a(rf_filter_coeff62_a), 
    .rf_filter_coeff62_b(rf_filter_coeff62_b), 
    .rf_filter_coeff63_a(rf_filter_coeff63_a), 
    .rf_filter_coeff63_b(rf_filter_coeff63_b), 
    .rf_filter_coeff64_a(rf_filter_coeff64_a), 
    .rf_filter_coeff64_b(rf_filter_coeff64_b), 
    .rf_filter_coeff65_a(rf_filter_coeff65_a), 
    .rf_filter_coeff65_b(rf_filter_coeff65_b), 
    .rf_filter_coeff66_a(rf_filter_coeff66_a), 
    .rf_filter_coeff66_b(rf_filter_coeff66_b), 
    .rf_filter_coeff67_a(rf_filter_coeff67_a), 
    .rf_filter_coeff67_b(rf_filter_coeff67_b), 
    .rf_filter_coeff68_a(rf_filter_coeff68_a), 
    .rf_filter_coeff68_b(rf_filter_coeff68_b), 
    .rf_filter_coeff69_a(rf_filter_coeff69_a), 
    .rf_filter_coeff69_b(rf_filter_coeff69_b), 
    .rf_filter_coeff70_a(rf_filter_coeff70_a), 
    .rf_filter_coeff70_b(rf_filter_coeff70_b), 
    .rf_filter_coeff71_a(rf_filter_coeff71_a), 
    .rf_filter_coeff71_b(rf_filter_coeff71_b), 
    .rf_filter_coeff72_a(rf_filter_coeff72_a), 
    .rf_filter_coeff72_b(rf_filter_coeff72_b), 
    .rf_filter_coeff73_a(rf_filter_coeff73_a), 
    .rf_filter_coeff73_b(rf_filter_coeff73_b), 
    .rf_filter_coeff74_a(rf_filter_coeff74_a), 
    .rf_filter_coeff74_b(rf_filter_coeff74_b), 
    .rf_filter_coeff75_a(rf_filter_coeff75_a), 
    .rf_filter_coeff75_b(rf_filter_coeff75_b), 
    .rf_filter_coeff76_a(rf_filter_coeff76_a), 
    .rf_filter_coeff76_b(rf_filter_coeff76_b), 
    .rf_filter_coeff77_a(rf_filter_coeff77_a), 
    .rf_filter_coeff77_b(rf_filter_coeff77_b), 
    .rf_filter_coeff78_a(rf_filter_coeff78_a), 
    .rf_filter_coeff78_b(rf_filter_coeff78_b), 
    .rf_filter_coeff79_a(rf_filter_coeff79_a), 
    .rf_filter_coeff79_b(rf_filter_coeff79_b), 
    .rf_filter_coeff80_a(rf_filter_coeff80_a), 
    .rf_filter_coeff80_b(rf_filter_coeff80_b), 
    .rf_filter_coeff81_a(rf_filter_coeff81_a), 
    .rf_filter_coeff81_b(rf_filter_coeff81_b), 
    .rf_filter_coeff82_a(rf_filter_coeff82_a), 
    .rf_filter_coeff82_b(rf_filter_coeff82_b), 
    .rf_filter_coeff83_a(rf_filter_coeff83_a), 
    .rf_filter_coeff83_b(rf_filter_coeff83_b), 
    .rf_filter_coeff84_a(rf_filter_coeff84_a), 
    .rf_filter_coeff84_b(rf_filter_coeff84_b), 
    .rf_filter_coeff85_a(rf_filter_coeff85_a), 
    .rf_filter_coeff85_b(rf_filter_coeff85_b), 
    .rf_filter_coeff86_a(rf_filter_coeff86_a), 
    .rf_filter_coeff86_b(rf_filter_coeff86_b), 
    .rf_filter_coeff87_a(rf_filter_coeff87_a), 
    .rf_filter_coeff87_b(rf_filter_coeff87_b), 
    .rf_filter_coeff88_a(rf_filter_coeff88_a), 
    .rf_filter_coeff88_b(rf_filter_coeff88_b), 
    .rf_filter_coeff89_a(rf_filter_coeff89_a), 
    .rf_filter_coeff89_b(rf_filter_coeff89_b), 
    .rf_filter_coeff90_a(rf_filter_coeff90_a), 
    .rf_filter_coeff90_b(rf_filter_coeff90_b), 
    .rf_filter_coeff91_a(rf_filter_coeff91_a), 
    .rf_filter_coeff91_b(rf_filter_coeff91_b), 
    .rf_filter_coeff92_a(rf_filter_coeff92_a), 
    .rf_filter_coeff92_b(rf_filter_coeff92_b), 
    .rf_filter_coeff93_a(rf_filter_coeff93_a), 
    .rf_filter_coeff93_b(rf_filter_coeff93_b), 
    .rf_filter_coeff94_a(rf_filter_coeff94_a), 
    .rf_filter_coeff94_b(rf_filter_coeff94_b), 
    .rf_filter_coeff95_a(rf_filter_coeff95_a), 
    .rf_filter_coeff95_b(rf_filter_coeff95_b), 
    .rf_filter_coeff96_a(rf_filter_coeff96_a), 
    .rf_filter_coeff96_b(rf_filter_coeff96_b), 
    .rf_filter_coeff97_a(rf_filter_coeff97_a), 
    .rf_filter_coeff97_b(rf_filter_coeff97_b), 
    .rf_filter_coeff98_a(rf_filter_coeff98_a), 
    .rf_filter_coeff98_b(rf_filter_coeff98_b), 
    .rf_filter_coeff99_a(rf_filter_coeff99_a), 
    .rf_filter_coeff99_b(rf_filter_coeff99_b), 
    .rf_filter_coeff100_a(rf_filter_coeff100_a), 
    .rf_filter_coeff100_b(rf_filter_coeff100_b), 
    .rf_filter_coeff101_a(rf_filter_coeff101_a), 
    .rf_filter_coeff101_b(rf_filter_coeff101_b), 
    .rf_filter_coeff102_a(rf_filter_coeff102_a), 
    .rf_filter_coeff102_b(rf_filter_coeff102_b), 
    .rf_filter_coeff103_a(rf_filter_coeff103_a), 
    .rf_filter_coeff103_b(rf_filter_coeff103_b), 
    .rf_filter_coeff104_a(rf_filter_coeff104_a), 
    .rf_filter_coeff104_b(rf_filter_coeff104_b), 
    .rf_filter_coeff105_a(rf_filter_coeff105_a), 
    .rf_filter_coeff105_b(rf_filter_coeff105_b), 
    .rf_filter_coeff106_a(rf_filter_coeff106_a), 
    .rf_filter_coeff106_b(rf_filter_coeff106_b), 
    .rf_filter_coeff107_a(rf_filter_coeff107_a), 
    .rf_filter_coeff107_b(rf_filter_coeff107_b), 
    .rf_filter_coeff108_a(rf_filter_coeff108_a), 
    .rf_filter_coeff108_b(rf_filter_coeff108_b), 
    .rf_filter_coeff109_a(rf_filter_coeff109_a), 
    .rf_filter_coeff109_b(rf_filter_coeff109_b), 
    .rf_filter_coeff110_a(rf_filter_coeff110_a), 
    .rf_filter_coeff110_b(rf_filter_coeff110_b), 
    .rf_filter_coeff111_a(rf_filter_coeff111_a), 
    .rf_filter_coeff111_b(rf_filter_coeff111_b), 
    .rf_filter_coeff112_a(rf_filter_coeff112_a), 
    .rf_filter_coeff112_b(rf_filter_coeff112_b), 
    .rf_filter_coeff113_a(rf_filter_coeff113_a), 
    .rf_filter_coeff113_b(rf_filter_coeff113_b), 
    .rf_filter_coeff114_a(rf_filter_coeff114_a), 
    .rf_filter_coeff114_b(rf_filter_coeff114_b), 
    .rf_filter_coeff115_a(rf_filter_coeff115_a), 
    .rf_filter_coeff115_b(rf_filter_coeff115_b), 
    .rf_filter_coeff116_a(rf_filter_coeff116_a), 
    .rf_filter_coeff116_b(rf_filter_coeff116_b), 
    .rf_filter_coeff117_a(rf_filter_coeff117_a), 
    .rf_filter_coeff117_b(rf_filter_coeff117_b), 
    .rf_filter_coeff118_a(rf_filter_coeff118_a), 
    .rf_filter_coeff118_b(rf_filter_coeff118_b), 
    .rf_filter_coeff119_a(rf_filter_coeff119_a), 
    .rf_filter_coeff119_b(rf_filter_coeff119_b), 
    .rf_filter_coeff120_a(rf_filter_coeff120_a), 
    .rf_filter_coeff120_b(rf_filter_coeff120_b), 
    .rf_filter_coeff121_a(rf_filter_coeff121_a), 
    .rf_filter_coeff121_b(rf_filter_coeff121_b), 
    .rf_filter_coeff122_a(rf_filter_coeff122_a), 
    .rf_filter_coeff122_b(rf_filter_coeff122_b), 
    .rf_filter_coeff123_a(rf_filter_coeff123_a), 
    .rf_filter_coeff123_b(rf_filter_coeff123_b), 
    .rf_filter_coeff124_a(rf_filter_coeff124_a), 
    .rf_filter_coeff124_b(rf_filter_coeff124_b), 
    .rf_filter_coeff125_a(rf_filter_coeff125_a), 
    .rf_filter_coeff125_b(rf_filter_coeff125_b), 
    .rf_filter_coeff126_a(rf_filter_coeff126_a), 
    .rf_filter_coeff126_b(rf_filter_coeff126_b), 
    .rf_filter_coeff127_a(rf_filter_coeff127_a), 
    .rf_filter_coeff127_b(rf_filter_coeff127_b), 
    .rf_filter_coeff128_a(rf_filter_coeff128_a), 
    .rf_filter_coeff128_b(rf_filter_coeff128_b), 
    .rf_filter_coeff129_a(rf_filter_coeff129_a), 
    .rf_filter_coeff129_b(rf_filter_coeff129_b), 
    .rf_filter_coeff130_a(rf_filter_coeff130_a), 
    .rf_filter_coeff130_b(rf_filter_coeff130_b), 
    .rf_filter_coeff131_a(rf_filter_coeff131_a), 
    .rf_filter_coeff131_b(rf_filter_coeff131_b), 
    .rf_filter_coeff132_a(rf_filter_coeff132_a), 
    .rf_filter_coeff132_b(rf_filter_coeff132_b), 
    .rf_filter_coeff133_a(rf_filter_coeff133_a), 
    .rf_filter_coeff133_b(rf_filter_coeff133_b), 
    .rf_filter_coeff134_a(rf_filter_coeff134_a), 
    .rf_filter_coeff134_b(rf_filter_coeff134_b), 
    .rf_filter_coeff135_a(rf_filter_coeff135_a), 
    .rf_filter_coeff135_b(rf_filter_coeff135_b), 
    .rf_filter_coeff136_a(rf_filter_coeff136_a), 
    .rf_filter_coeff136_b(rf_filter_coeff136_b), 
    .rf_filter_coeff137_a(rf_filter_coeff137_a), 
    .rf_filter_coeff137_b(rf_filter_coeff137_b), 
    .rf_filter_coeff138_a(rf_filter_coeff138_a), 
    .rf_filter_coeff138_b(rf_filter_coeff138_b), 
    .rf_filter_coeff139_a(rf_filter_coeff139_a), 
    .rf_filter_coeff139_b(rf_filter_coeff139_b), 
    .rf_filter_coeff140_a(rf_filter_coeff140_a), 
    .rf_filter_coeff140_b(rf_filter_coeff140_b), 
    .rf_filter_coeff141_a(rf_filter_coeff141_a), 
    .rf_filter_coeff141_b(rf_filter_coeff141_b), 
    .rf_filter_coeff142_a(rf_filter_coeff142_a), 
    .rf_filter_coeff142_b(rf_filter_coeff142_b), 
    .rf_filter_coeff143_a(rf_filter_coeff143_a), 
    .rf_filter_coeff143_b(rf_filter_coeff143_b), 
    .rf_filter_coeff144_a(rf_filter_coeff144_a), 
    .rf_filter_coeff144_b(rf_filter_coeff144_b), 
    .rf_filter_coeff145_a(rf_filter_coeff145_a), 
    .rf_filter_coeff145_b(rf_filter_coeff145_b), 
    .rf_filter_coeff146_a(rf_filter_coeff146_a), 
    .rf_filter_coeff146_b(rf_filter_coeff146_b), 
    .rf_filter_coeff147_a(rf_filter_coeff147_a), 
    .rf_filter_coeff147_b(rf_filter_coeff147_b), 
    .rf_filter_coeff148_a(rf_filter_coeff148_a), 
    .rf_filter_coeff148_b(rf_filter_coeff148_b), 
    .rf_filter_coeff149_a(rf_filter_coeff149_a), 
    .rf_filter_coeff149_b(rf_filter_coeff149_b), 
    .rf_filter_coeff150_a(rf_filter_coeff150_a), 
    .rf_filter_coeff150_b(rf_filter_coeff150_b), 
    .rf_filter_coeff151_a(rf_filter_coeff151_a), 
    .rf_filter_coeff151_b(rf_filter_coeff151_b), 
    .rf_filter_coeff152_a(rf_filter_coeff152_a), 
    .rf_filter_coeff152_b(rf_filter_coeff152_b), 
    .rf_filter_coeff153_a(rf_filter_coeff153_a), 
    .rf_filter_coeff153_b(rf_filter_coeff153_b), 
    .rf_filter_coeff154_a(rf_filter_coeff154_a), 
    .rf_filter_coeff154_b(rf_filter_coeff154_b), 
    .rf_filter_coeff155_a(rf_filter_coeff155_a), 
    .rf_filter_coeff155_b(rf_filter_coeff155_b), 
    .rf_filter_coeff156_a(rf_filter_coeff156_a), 
    .rf_filter_coeff156_b(rf_filter_coeff156_b), 
    .rf_filter_coeff157_a(rf_filter_coeff157_a), 
    .rf_filter_coeff157_b(rf_filter_coeff157_b), 
    .rf_filter_coeff158_a(rf_filter_coeff158_a), 
    .rf_filter_coeff158_b(rf_filter_coeff158_b), 
    .rf_filter_coeff159_a(rf_filter_coeff159_a), 
    .rf_filter_coeff159_b(rf_filter_coeff159_b), 
    .rf_filter_coeff160_a(rf_filter_coeff160_a), 
    .rf_filter_coeff160_b(rf_filter_coeff160_b), 
    .rf_filter_coeff161_a(rf_filter_coeff161_a), 
    .rf_filter_coeff161_b(rf_filter_coeff161_b), 
    .rf_filter_coeff162_a(rf_filter_coeff162_a), 
    .rf_filter_coeff162_b(rf_filter_coeff162_b), 
    .rf_filter_coeff163_a(rf_filter_coeff163_a), 
    .rf_filter_coeff163_b(rf_filter_coeff163_b), 
    .rf_filter_coeff164_a(rf_filter_coeff164_a), 
    .rf_filter_coeff164_b(rf_filter_coeff164_b), 
    .rf_filter_coeff165_a(rf_filter_coeff165_a), 
    .rf_filter_coeff165_b(rf_filter_coeff165_b), 
    .rf_filter_coeff166_a(rf_filter_coeff166_a), 
    .rf_filter_coeff166_b(rf_filter_coeff166_b), 
    .rf_filter_coeff167_a(rf_filter_coeff167_a), 
    .rf_filter_coeff167_b(rf_filter_coeff167_b), 
    .rf_filter_coeff168_a(rf_filter_coeff168_a), 
    .rf_filter_coeff168_b(rf_filter_coeff168_b), 
    .rf_filter_coeff169_a(rf_filter_coeff169_a), 
    .rf_filter_coeff169_b(rf_filter_coeff169_b), 
    .rf_filter_coeff170_a(rf_filter_coeff170_a), 
    .rf_filter_coeff170_b(rf_filter_coeff170_b), 
    .rf_filter_coeff171_a(rf_filter_coeff171_a), 
    .rf_filter_coeff171_b(rf_filter_coeff171_b), 
    .rf_filter_coeff172_a(rf_filter_coeff172_a), 
    .rf_filter_coeff172_b(rf_filter_coeff172_b), 
    .rf_filter_coeff173_a(rf_filter_coeff173_a), 
    .rf_filter_coeff173_b(rf_filter_coeff173_b), 
    .rf_filter_coeff174_a(rf_filter_coeff174_a), 
    .rf_filter_coeff174_b(rf_filter_coeff174_b), 
    .rf_filter_coeff175_a(rf_filter_coeff175_a), 
    .rf_filter_coeff175_b(rf_filter_coeff175_b), 
    .rf_filter_coeff176_a(rf_filter_coeff176_a), 
    .rf_filter_coeff176_b(rf_filter_coeff176_b), 
    .rf_filter_coeff177_a(rf_filter_coeff177_a), 
    .rf_filter_coeff177_b(rf_filter_coeff177_b), 
    .rf_filter_coeff178_a(rf_filter_coeff178_a), 
    .rf_filter_coeff178_b(rf_filter_coeff178_b), 
    .rf_filter_coeff179_a(rf_filter_coeff179_a), 
    .rf_filter_coeff179_b(rf_filter_coeff179_b), 
    .rf_filter_coeff180_a(rf_filter_coeff180_a), 
    .rf_filter_coeff180_b(rf_filter_coeff180_b), 
    .rf_filter_coeff181_a(rf_filter_coeff181_a), 
    .rf_filter_coeff181_b(rf_filter_coeff181_b), 
    .rf_filter_coeff182_a(rf_filter_coeff182_a), 
    .rf_filter_coeff182_b(rf_filter_coeff182_b), 
    .rf_filter_coeff183_a(rf_filter_coeff183_a), 
    .rf_filter_coeff183_b(rf_filter_coeff183_b), 
    .rf_filter_coeff184_a(rf_filter_coeff184_a), 
    .rf_filter_coeff184_b(rf_filter_coeff184_b), 
    .rf_filter_coeff185_a(rf_filter_coeff185_a), 
    .rf_filter_coeff185_b(rf_filter_coeff185_b), 
    .rf_filter_coeff186_a(rf_filter_coeff186_a), 
    .rf_filter_coeff186_b(rf_filter_coeff186_b), 
    .rf_filter_coeff187_a(rf_filter_coeff187_a), 
    .rf_filter_coeff187_b(rf_filter_coeff187_b), 
    .rf_filter_coeff188_a(rf_filter_coeff188_a), 
    .rf_filter_coeff188_b(rf_filter_coeff188_b), 
    .rf_filter_coeff189_a(rf_filter_coeff189_a), 
    .rf_filter_coeff189_b(rf_filter_coeff189_b), 
    .rf_filter_coeff190_a(rf_filter_coeff190_a), 
    .rf_filter_coeff190_b(rf_filter_coeff190_b), 
    .rf_filter_coeff191_a(rf_filter_coeff191_a), 
    .rf_filter_coeff191_b(rf_filter_coeff191_b), 
    .rf_filter_coeff192_a(rf_filter_coeff192_a), 
    .rf_filter_coeff192_b(rf_filter_coeff192_b), 
    .rf_filter_coeff193_a(rf_filter_coeff193_a), 
    .rf_filter_coeff193_b(rf_filter_coeff193_b), 
    .rf_filter_coeff194_a(rf_filter_coeff194_a), 
    .rf_filter_coeff194_b(rf_filter_coeff194_b), 
    .rf_filter_coeff195_a(rf_filter_coeff195_a), 
    .rf_filter_coeff195_b(rf_filter_coeff195_b), 
    .rf_filter_coeff196_a(rf_filter_coeff196_a), 
    .rf_filter_coeff196_b(rf_filter_coeff196_b), 
    .rf_filter_coeff197_a(rf_filter_coeff197_a), 
    .rf_filter_coeff197_b(rf_filter_coeff197_b), 
    .rf_filter_coeff198_a(rf_filter_coeff198_a), 
    .rf_filter_coeff198_b(rf_filter_coeff198_b), 
    .rf_filter_coeff199_a(rf_filter_coeff199_a), 
    .rf_filter_coeff199_b(rf_filter_coeff199_b), 
    .rf_filter_coeff200_a(rf_filter_coeff200_a), 
    .rf_filter_coeff200_b(rf_filter_coeff200_b), 
    .rf_filter_coeff201_a(rf_filter_coeff201_a), 
    .rf_filter_coeff201_b(rf_filter_coeff201_b), 
    .rf_filter_coeff202_a(rf_filter_coeff202_a), 
    .rf_filter_coeff202_b(rf_filter_coeff202_b), 
    .rf_filter_coeff203_a(rf_filter_coeff203_a), 
    .rf_filter_coeff203_b(rf_filter_coeff203_b), 
    .rf_filter_coeff204_a(rf_filter_coeff204_a), 
    .rf_filter_coeff204_b(rf_filter_coeff204_b), 
    .rf_filter_coeff205_a(rf_filter_coeff205_a), 
    .rf_filter_coeff205_b(rf_filter_coeff205_b), 
    .rf_filter_coeff206_a(rf_filter_coeff206_a), 
    .rf_filter_coeff206_b(rf_filter_coeff206_b), 
    .rf_filter_coeff207_a(rf_filter_coeff207_a), 
    .rf_filter_coeff207_b(rf_filter_coeff207_b), 
    .rf_filter_coeff208_a(rf_filter_coeff208_a), 
    .rf_filter_coeff208_b(rf_filter_coeff208_b), 
    .rf_filter_coeff209_a(rf_filter_coeff209_a), 
    .rf_filter_coeff209_b(rf_filter_coeff209_b), 
    .rf_filter_coeff210_a(rf_filter_coeff210_a), 
    .rf_filter_coeff210_b(rf_filter_coeff210_b), 
    .rf_filter_coeff211_a(rf_filter_coeff211_a), 
    .rf_filter_coeff211_b(rf_filter_coeff211_b), 
    .rf_filter_coeff212_a(rf_filter_coeff212_a), 
    .rf_filter_coeff212_b(rf_filter_coeff212_b), 
    .rf_filter_coeff213_a(rf_filter_coeff213_a), 
    .rf_filter_coeff213_b(rf_filter_coeff213_b), 
    .rf_filter_coeff214_a(rf_filter_coeff214_a), 
    .rf_filter_coeff214_b(rf_filter_coeff214_b), 
    .rf_filter_coeff215_a(rf_filter_coeff215_a), 
    .rf_filter_coeff215_b(rf_filter_coeff215_b), 
    .rf_filter_coeff216_a(rf_filter_coeff216_a), 
    .rf_filter_coeff216_b(rf_filter_coeff216_b), 
    .rf_filter_coeff217_a(rf_filter_coeff217_a), 
    .rf_filter_coeff217_b(rf_filter_coeff217_b), 
    .rf_filter_coeff218_a(rf_filter_coeff218_a), 
    .rf_filter_coeff218_b(rf_filter_coeff218_b), 
    .rf_filter_coeff219_a(rf_filter_coeff219_a), 
    .rf_filter_coeff219_b(rf_filter_coeff219_b), 
    .rf_filter_coeff220_a(rf_filter_coeff220_a), 
    .rf_filter_coeff220_b(rf_filter_coeff220_b), 
    .rf_filter_coeff221_a(rf_filter_coeff221_a), 
    .rf_filter_coeff221_b(rf_filter_coeff221_b), 
    .rf_filter_coeff222_a(rf_filter_coeff222_a), 
    .rf_filter_coeff222_b(rf_filter_coeff222_b), 
    .rf_filter_coeff223_a(rf_filter_coeff223_a), 
    .rf_filter_coeff223_b(rf_filter_coeff223_b), 
    .rf_filter_coeff224_a(rf_filter_coeff224_a), 
    .rf_filter_coeff224_b(rf_filter_coeff224_b), 
    .rf_filter_coeff225_a(rf_filter_coeff225_a), 
    .rf_filter_coeff225_b(rf_filter_coeff225_b), 
    .rf_filter_coeff226_a(rf_filter_coeff226_a), 
    .rf_filter_coeff226_b(rf_filter_coeff226_b), 
    .rf_filter_coeff227_a(rf_filter_coeff227_a), 
    .rf_filter_coeff227_b(rf_filter_coeff227_b), 
    .rf_filter_coeff228_a(rf_filter_coeff228_a), 
    .rf_filter_coeff228_b(rf_filter_coeff228_b), 
    .rf_filter_coeff229_a(rf_filter_coeff229_a), 
    .rf_filter_coeff229_b(rf_filter_coeff229_b), 
    .rf_filter_coeff230_a(rf_filter_coeff230_a), 
    .rf_filter_coeff230_b(rf_filter_coeff230_b), 
    .rf_filter_coeff231_a(rf_filter_coeff231_a), 
    .rf_filter_coeff231_b(rf_filter_coeff231_b), 
    .rf_filter_coeff232_a(rf_filter_coeff232_a), 
    .rf_filter_coeff232_b(rf_filter_coeff232_b), 
    .rf_filter_coeff233_a(rf_filter_coeff233_a), 
    .rf_filter_coeff233_b(rf_filter_coeff233_b), 
    .rf_filter_coeff234_a(rf_filter_coeff234_a), 
    .rf_filter_coeff234_b(rf_filter_coeff234_b), 
    .rf_filter_coeff235_a(rf_filter_coeff235_a), 
    .rf_filter_coeff235_b(rf_filter_coeff235_b), 
    .rf_filter_coeff236_a(rf_filter_coeff236_a), 
    .rf_filter_coeff236_b(rf_filter_coeff236_b), 
    .rf_filter_coeff237_a(rf_filter_coeff237_a), 
    .rf_filter_coeff237_b(rf_filter_coeff237_b), 
    .rf_filter_coeff238_a(rf_filter_coeff238_a), 
    .rf_filter_coeff238_b(rf_filter_coeff238_b), 
    .rf_filter_coeff239_a(rf_filter_coeff239_a), 
    .rf_filter_coeff239_b(rf_filter_coeff239_b), 
    .rf_filter_coeff240_a(rf_filter_coeff240_a), 
    .rf_filter_coeff240_b(rf_filter_coeff240_b), 
    .rf_filter_coeff241_a(rf_filter_coeff241_a), 
    .rf_filter_coeff241_b(rf_filter_coeff241_b), 
    .rf_filter_coeff242_a(rf_filter_coeff242_a), 
    .rf_filter_coeff242_b(rf_filter_coeff242_b), 
    .rf_filter_coeff243_a(rf_filter_coeff243_a), 
    .rf_filter_coeff243_b(rf_filter_coeff243_b), 
    .rf_filter_coeff244_a(rf_filter_coeff244_a), 
    .rf_filter_coeff244_b(rf_filter_coeff244_b), 
    .rf_filter_coeff245_a(rf_filter_coeff245_a), 
    .rf_filter_coeff245_b(rf_filter_coeff245_b), 
    .rf_filter_coeff246_a(rf_filter_coeff246_a), 
    .rf_filter_coeff246_b(rf_filter_coeff246_b), 
    .rf_filter_coeff247_a(rf_filter_coeff247_a), 
    .rf_filter_coeff247_b(rf_filter_coeff247_b), 
    .rf_filter_coeff248_a(rf_filter_coeff248_a), 
    .rf_filter_coeff248_b(rf_filter_coeff248_b), 
    .rf_filter_coeff249_a(rf_filter_coeff249_a), 
    .rf_filter_coeff249_b(rf_filter_coeff249_b), 
    .rf_filter_coeff250_a(rf_filter_coeff250_a), 
    .rf_filter_coeff250_b(rf_filter_coeff250_b), 
    .rf_filter_coeff251_a(rf_filter_coeff251_a), 
    .rf_filter_coeff251_b(rf_filter_coeff251_b), 
    .rf_filter_coeff252_a(rf_filter_coeff252_a), 
    .rf_filter_coeff252_b(rf_filter_coeff252_b), 
    .rf_filter_coeff253_a(rf_filter_coeff253_a), 
    .rf_filter_coeff253_b(rf_filter_coeff253_b), 
    .rf_filter_coeff254_a(rf_filter_coeff254_a), 
    .rf_filter_coeff254_b(rf_filter_coeff254_b), 
    .rf_filter_coeff255_a(rf_filter_coeff255_a), 
    .rf_filter_coeff255_b(rf_filter_coeff255_b), 
    .rf_filter_coeff256_a(rf_filter_coeff256_a), 
    .rf_filter_coeff256_b(rf_filter_coeff256_b), 
    .rf_filter_coeff257_a(rf_filter_coeff257_a), 
    .rf_filter_coeff257_b(rf_filter_coeff257_b), 
    .rf_filter_coeff258_a(rf_filter_coeff258_a), 
    .rf_filter_coeff258_b(rf_filter_coeff258_b), 
    .rf_filter_coeff259_a(rf_filter_coeff259_a), 
    .rf_filter_coeff259_b(rf_filter_coeff259_b), 
    .rf_filter_coeff260_a(rf_filter_coeff260_a), 
    .rf_filter_coeff260_b(rf_filter_coeff260_b), 
    .rf_filter_coeff261_a(rf_filter_coeff261_a), 
    .rf_filter_coeff261_b(rf_filter_coeff261_b), 
    .rf_filter_coeff262_a(rf_filter_coeff262_a), 
    .rf_filter_coeff262_b(rf_filter_coeff262_b), 
    .rf_filter_coeff263_a(rf_filter_coeff263_a), 
    .rf_filter_coeff263_b(rf_filter_coeff263_b), 
    .rf_filter_coeff264_a(rf_filter_coeff264_a), 
    .rf_filter_coeff264_b(rf_filter_coeff264_b), 
    .rf_filter_coeff265_a(rf_filter_coeff265_a), 
    .rf_filter_coeff265_b(rf_filter_coeff265_b), 
    .rf_filter_coeff266_a(rf_filter_coeff266_a), 
    .rf_filter_coeff266_b(rf_filter_coeff266_b), 
    .rf_filter_coeff267_a(rf_filter_coeff267_a), 
    .rf_filter_coeff267_b(rf_filter_coeff267_b), 
    .rf_filter_coeff268_a(rf_filter_coeff268_a), 
    .rf_filter_coeff268_b(rf_filter_coeff268_b), 
    .rf_filter_coeff269_a(rf_filter_coeff269_a), 
    .rf_filter_coeff269_b(rf_filter_coeff269_b), 
    .rf_filter_coeff270_a(rf_filter_coeff270_a), 
    .rf_filter_coeff270_b(rf_filter_coeff270_b), 
    .rf_filter_coeff271_a(rf_filter_coeff271_a), 
    .rf_filter_coeff271_b(rf_filter_coeff271_b), 
    .rf_filter_coeff272_a(rf_filter_coeff272_a), 
    .rf_filter_coeff272_b(rf_filter_coeff272_b), 
    .rf_filter_coeff273_a(rf_filter_coeff273_a), 
    .rf_filter_coeff273_b(rf_filter_coeff273_b), 
    .rf_filter_coeff274_a(rf_filter_coeff274_a), 
    .rf_filter_coeff274_b(rf_filter_coeff274_b), 
    .rf_filter_coeff275_a(rf_filter_coeff275_a), 
    .rf_filter_coeff275_b(rf_filter_coeff275_b), 
    .rf_filter_coeff276_a(rf_filter_coeff276_a), 
    .rf_filter_coeff276_b(rf_filter_coeff276_b), 
    .rf_filter_coeff277_a(rf_filter_coeff277_a), 
    .rf_filter_coeff277_b(rf_filter_coeff277_b), 
    .rf_filter_coeff278_a(rf_filter_coeff278_a), 
    .rf_filter_coeff278_b(rf_filter_coeff278_b), 
    .rf_filter_coeff279_a(rf_filter_coeff279_a), 
    .rf_filter_coeff279_b(rf_filter_coeff279_b), 
    .rf_filter_coeff280_a(rf_filter_coeff280_a), 
    .rf_filter_coeff280_b(rf_filter_coeff280_b), 
    .rf_filter_coeff281_a(rf_filter_coeff281_a), 
    .rf_filter_coeff281_b(rf_filter_coeff281_b), 
    .rf_filter_coeff282_a(rf_filter_coeff282_a), 
    .rf_filter_coeff282_b(rf_filter_coeff282_b), 
    .rf_filter_coeff283_a(rf_filter_coeff283_a), 
    .rf_filter_coeff283_b(rf_filter_coeff283_b), 
    .rf_filter_coeff284_a(rf_filter_coeff284_a), 
    .rf_filter_coeff284_b(rf_filter_coeff284_b), 
    .rf_filter_coeff285_a(rf_filter_coeff285_a), 
    .rf_filter_coeff285_b(rf_filter_coeff285_b), 
    .rf_filter_coeff286_a(rf_filter_coeff286_a), 
    .rf_filter_coeff286_b(rf_filter_coeff286_b), 
    .rf_filter_coeff287_a(rf_filter_coeff287_a), 
    .rf_filter_coeff287_b(rf_filter_coeff287_b), 
    .rf_filter_coeff288_a(rf_filter_coeff288_a), 
    .rf_filter_coeff288_b(rf_filter_coeff288_b), 
    .rf_filter_coeff289_a(rf_filter_coeff289_a), 
    .rf_filter_coeff289_b(rf_filter_coeff289_b), 
    .rf_filter_coeff290_a(rf_filter_coeff290_a), 
    .rf_filter_coeff290_b(rf_filter_coeff290_b), 
    .rf_filter_coeff291_a(rf_filter_coeff291_a), 
    .rf_filter_coeff291_b(rf_filter_coeff291_b), 
    .rf_filter_coeff292_a(rf_filter_coeff292_a), 
    .rf_filter_coeff292_b(rf_filter_coeff292_b), 
    .rf_filter_coeff293_a(rf_filter_coeff293_a), 
    .rf_filter_coeff293_b(rf_filter_coeff293_b), 
    .rf_filter_coeff294_a(rf_filter_coeff294_a), 
    .rf_filter_coeff294_b(rf_filter_coeff294_b), 
    .rf_filter_coeff295_a(rf_filter_coeff295_a), 
    .rf_filter_coeff295_b(rf_filter_coeff295_b), 
    .rf_filter_coeff296_a(rf_filter_coeff296_a), 
    .rf_filter_coeff296_b(rf_filter_coeff296_b), 
    .rf_filter_coeff297_a(rf_filter_coeff297_a), 
    .rf_filter_coeff297_b(rf_filter_coeff297_b), 
    .rf_filter_coeff298_a(rf_filter_coeff298_a), 
    .rf_filter_coeff298_b(rf_filter_coeff298_b), 
    .rf_filter_coeff299_a(rf_filter_coeff299_a), 
    .rf_filter_coeff299_b(rf_filter_coeff299_b), 
    .rf_filter_coeff300_a(rf_filter_coeff300_a), 
    .rf_filter_coeff300_b(rf_filter_coeff300_b), 
    .rf_filter_coeff301_a(rf_filter_coeff301_a), 
    .rf_filter_coeff301_b(rf_filter_coeff301_b), 
    .rf_filter_coeff302_a(rf_filter_coeff302_a), 
    .rf_filter_coeff302_b(rf_filter_coeff302_b), 
    .rf_filter_coeff303_a(rf_filter_coeff303_a), 
    .rf_filter_coeff303_b(rf_filter_coeff303_b), 
    .rf_filter_coeff304_a(rf_filter_coeff304_a), 
    .rf_filter_coeff304_b(rf_filter_coeff304_b), 
    .rf_filter_coeff305_a(rf_filter_coeff305_a), 
    .rf_filter_coeff305_b(rf_filter_coeff305_b), 
    .rf_filter_coeff306_a(rf_filter_coeff306_a), 
    .rf_filter_coeff306_b(rf_filter_coeff306_b), 
    .rf_filter_coeff307_a(rf_filter_coeff307_a), 
    .rf_filter_coeff307_b(rf_filter_coeff307_b), 
    .rf_filter_coeff308_a(rf_filter_coeff308_a), 
    .rf_filter_coeff308_b(rf_filter_coeff308_b), 
    .rf_filter_coeff309_a(rf_filter_coeff309_a), 
    .rf_filter_coeff309_b(rf_filter_coeff309_b), 
    .rf_filter_coeff310_a(rf_filter_coeff310_a), 
    .rf_filter_coeff310_b(rf_filter_coeff310_b), 
    .rf_filter_coeff311_a(rf_filter_coeff311_a), 
    .rf_filter_coeff311_b(rf_filter_coeff311_b), 
    .rf_filter_coeff312_a(rf_filter_coeff312_a), 
    .rf_filter_coeff312_b(rf_filter_coeff312_b), 
    .rf_filter_coeff313_a(rf_filter_coeff313_a), 
    .rf_filter_coeff313_b(rf_filter_coeff313_b), 
    .rf_filter_coeff314_a(rf_filter_coeff314_a), 
    .rf_filter_coeff314_b(rf_filter_coeff314_b), 
    .rf_filter_coeff315_a(rf_filter_coeff315_a), 
    .rf_filter_coeff315_b(rf_filter_coeff315_b), 
    .rf_filter_coeff316_a(rf_filter_coeff316_a), 
    .rf_filter_coeff316_b(rf_filter_coeff316_b), 
    .rf_filter_coeff317_a(rf_filter_coeff317_a), 
    .rf_filter_coeff317_b(rf_filter_coeff317_b), 
    .rf_filter_coeff318_a(rf_filter_coeff318_a), 
    .rf_filter_coeff318_b(rf_filter_coeff318_b), 
    .rf_filter_coeff319_a(rf_filter_coeff319_a), 
    .rf_filter_coeff319_b(rf_filter_coeff319_b), 
    .rf_filter_coeff320_a(rf_filter_coeff320_a), 
    .rf_filter_coeff320_b(rf_filter_coeff320_b), 
    .rf_filter_coeff321_a(rf_filter_coeff321_a), 
    .rf_filter_coeff321_b(rf_filter_coeff321_b), 
    .rf_filter_coeff322_a(rf_filter_coeff322_a), 
    .rf_filter_coeff322_b(rf_filter_coeff322_b), 
    .rf_filter_coeff323_a(rf_filter_coeff323_a), 
    .rf_filter_coeff323_b(rf_filter_coeff323_b), 
    .rf_filter_coeff324_a(rf_filter_coeff324_a), 
    .rf_filter_coeff324_b(rf_filter_coeff324_b), 
    .rf_filter_coeff325_a(rf_filter_coeff325_a), 
    .rf_filter_coeff325_b(rf_filter_coeff325_b), 
    .rf_filter_coeff326_a(rf_filter_coeff326_a), 
    .rf_filter_coeff326_b(rf_filter_coeff326_b), 
    .rf_filter_coeff327_a(rf_filter_coeff327_a), 
    .rf_filter_coeff327_b(rf_filter_coeff327_b), 
    .rf_filter_coeff328_a(rf_filter_coeff328_a), 
    .rf_filter_coeff328_b(rf_filter_coeff328_b), 
    .rf_filter_coeff329_a(rf_filter_coeff329_a), 
    .rf_filter_coeff329_b(rf_filter_coeff329_b), 
    .rf_filter_coeff330_a(rf_filter_coeff330_a), 
    .rf_filter_coeff330_b(rf_filter_coeff330_b), 
    .rf_filter_coeff331_a(rf_filter_coeff331_a), 
    .rf_filter_coeff331_b(rf_filter_coeff331_b), 
    .rf_filter_coeff332_a(rf_filter_coeff332_a), 
    .rf_filter_coeff332_b(rf_filter_coeff332_b), 
    .rf_filter_coeff333_a(rf_filter_coeff333_a), 
    .rf_filter_coeff333_b(rf_filter_coeff333_b), 
    .rf_filter_coeff334_a(rf_filter_coeff334_a), 
    .rf_filter_coeff334_b(rf_filter_coeff334_b), 
    .rf_filter_coeff335_a(rf_filter_coeff335_a), 
    .rf_filter_coeff335_b(rf_filter_coeff335_b), 
    .rf_filter_coeff336_a(rf_filter_coeff336_a), 
    .rf_filter_coeff336_b(rf_filter_coeff336_b), 
    .rf_filter_coeff337_a(rf_filter_coeff337_a), 
    .rf_filter_coeff337_b(rf_filter_coeff337_b), 
    .rf_filter_coeff338_a(rf_filter_coeff338_a), 
    .rf_filter_coeff338_b(rf_filter_coeff338_b), 
    .rf_filter_coeff339_a(rf_filter_coeff339_a), 
    .rf_filter_coeff339_b(rf_filter_coeff339_b), 
    .rf_filter_coeff340_a(rf_filter_coeff340_a), 
    .rf_filter_coeff340_b(rf_filter_coeff340_b), 
    .rf_filter_coeff341_a(rf_filter_coeff341_a), 
    .rf_filter_coeff341_b(rf_filter_coeff341_b), 
    .rf_filter_coeff342_a(rf_filter_coeff342_a), 
    .rf_filter_coeff342_b(rf_filter_coeff342_b), 
    .rf_filter_coeff343_a(rf_filter_coeff343_a), 
    .rf_filter_coeff343_b(rf_filter_coeff343_b), 
    .rf_filter_coeff344_a(rf_filter_coeff344_a), 
    .rf_filter_coeff344_b(rf_filter_coeff344_b), 
    .rf_filter_coeff345_a(rf_filter_coeff345_a), 
    .rf_filter_coeff345_b(rf_filter_coeff345_b), 
    .rf_filter_coeff346_a(rf_filter_coeff346_a), 
    .rf_filter_coeff346_b(rf_filter_coeff346_b), 
    .rf_filter_coeff347_a(rf_filter_coeff347_a), 
    .rf_filter_coeff347_b(rf_filter_coeff347_b), 
    .rf_filter_coeff348_a(rf_filter_coeff348_a), 
    .rf_filter_coeff348_b(rf_filter_coeff348_b), 
    .rf_filter_coeff349_a(rf_filter_coeff349_a), 
    .rf_filter_coeff349_b(rf_filter_coeff349_b), 
    .rf_filter_coeff350_a(rf_filter_coeff350_a), 
    .rf_filter_coeff350_b(rf_filter_coeff350_b), 
    .rf_filter_coeff351_a(rf_filter_coeff351_a), 
    .rf_filter_coeff351_b(rf_filter_coeff351_b), 
    .rf_filter_coeff352_a(rf_filter_coeff352_a), 
    .rf_filter_coeff352_b(rf_filter_coeff352_b), 
    .rf_filter_coeff353_a(rf_filter_coeff353_a), 
    .rf_filter_coeff353_b(rf_filter_coeff353_b), 
    .rf_filter_coeff354_a(rf_filter_coeff354_a), 
    .rf_filter_coeff354_b(rf_filter_coeff354_b), 
    .rf_filter_coeff355_a(rf_filter_coeff355_a), 
    .rf_filter_coeff355_b(rf_filter_coeff355_b), 
    .rf_filter_coeff356_a(rf_filter_coeff356_a), 
    .rf_filter_coeff356_b(rf_filter_coeff356_b), 
    .rf_filter_coeff357_a(rf_filter_coeff357_a), 
    .rf_filter_coeff357_b(rf_filter_coeff357_b), 
    .rf_filter_coeff358_a(rf_filter_coeff358_a), 
    .rf_filter_coeff358_b(rf_filter_coeff358_b), 
    .rf_filter_coeff359_a(rf_filter_coeff359_a), 
    .rf_filter_coeff359_b(rf_filter_coeff359_b), 
    .rf_filter_coeff360_a(rf_filter_coeff360_a), 
    .rf_filter_coeff360_b(rf_filter_coeff360_b), 
    .rf_filter_coeff361_a(rf_filter_coeff361_a), 
    .rf_filter_coeff361_b(rf_filter_coeff361_b), 
    .rf_filter_coeff362_a(rf_filter_coeff362_a), 
    .rf_filter_coeff362_b(rf_filter_coeff362_b), 
    .rf_filter_coeff363_a(rf_filter_coeff363_a), 
    .rf_filter_coeff363_b(rf_filter_coeff363_b), 
    .rf_filter_coeff364_a(rf_filter_coeff364_a), 
    .rf_filter_coeff364_b(rf_filter_coeff364_b), 
    .rf_filter_coeff365_a(rf_filter_coeff365_a), 
    .rf_filter_coeff365_b(rf_filter_coeff365_b), 
    .rf_filter_coeff366_a(rf_filter_coeff366_a), 
    .rf_filter_coeff366_b(rf_filter_coeff366_b), 
    .rf_filter_coeff367_a(rf_filter_coeff367_a), 
    .rf_filter_coeff367_b(rf_filter_coeff367_b), 
    .rf_filter_coeff368_a(rf_filter_coeff368_a), 
    .rf_filter_coeff368_b(rf_filter_coeff368_b), 
    .rf_filter_coeff369_a(rf_filter_coeff369_a), 
    .rf_filter_coeff369_b(rf_filter_coeff369_b), 
    .rf_filter_coeff370_a(rf_filter_coeff370_a), 
    .rf_filter_coeff370_b(rf_filter_coeff370_b), 
    .rf_filter_coeff371_a(rf_filter_coeff371_a), 
    .rf_filter_coeff371_b(rf_filter_coeff371_b), 
    .rf_filter_coeff372_a(rf_filter_coeff372_a), 
    .rf_filter_coeff372_b(rf_filter_coeff372_b), 
    .rf_filter_coeff373_a(rf_filter_coeff373_a), 
    .rf_filter_coeff373_b(rf_filter_coeff373_b), 
    .rf_filter_coeff374_a(rf_filter_coeff374_a), 
    .rf_filter_coeff374_b(rf_filter_coeff374_b), 
    .rf_filter_coeff375_a(rf_filter_coeff375_a), 
    .rf_filter_coeff375_b(rf_filter_coeff375_b), 
    .rf_filter_coeff376_a(rf_filter_coeff376_a), 
    .rf_filter_coeff376_b(rf_filter_coeff376_b), 
    .rf_filter_coeff377_a(rf_filter_coeff377_a), 
    .rf_filter_coeff377_b(rf_filter_coeff377_b), 
    .rf_filter_coeff378_a(rf_filter_coeff378_a), 
    .rf_filter_coeff378_b(rf_filter_coeff378_b), 
    .rf_filter_coeff379_a(rf_filter_coeff379_a), 
    .rf_filter_coeff379_b(rf_filter_coeff379_b), 
    .rf_filter_coeff380_a(rf_filter_coeff380_a), 
    .rf_filter_coeff380_b(rf_filter_coeff380_b), 
    .rf_filter_coeff381_a(rf_filter_coeff381_a), 
    .rf_filter_coeff381_b(rf_filter_coeff381_b), 
    .rf_filter_coeff382_a(rf_filter_coeff382_a), 
    .rf_filter_coeff382_b(rf_filter_coeff382_b), 
    .rf_filter_coeff383_a(rf_filter_coeff383_a), 
    .rf_filter_coeff383_b(rf_filter_coeff383_b), 
    .rf_filter_coeff384_a(rf_filter_coeff384_a), 
    .rf_filter_coeff384_b(rf_filter_coeff384_b), 
    .rf_filter_coeff385_a(rf_filter_coeff385_a), 
    .rf_filter_coeff385_b(rf_filter_coeff385_b), 
    .rf_filter_coeff386_a(rf_filter_coeff386_a), 
    .rf_filter_coeff386_b(rf_filter_coeff386_b), 
    .rf_filter_coeff387_a(rf_filter_coeff387_a), 
    .rf_filter_coeff387_b(rf_filter_coeff387_b), 
    .rf_filter_coeff388_a(rf_filter_coeff388_a), 
    .rf_filter_coeff388_b(rf_filter_coeff388_b), 
    .rf_filter_coeff389_a(rf_filter_coeff389_a), 
    .rf_filter_coeff389_b(rf_filter_coeff389_b), 
    .rf_filter_coeff390_a(rf_filter_coeff390_a), 
    .rf_filter_coeff390_b(rf_filter_coeff390_b), 
    .rf_filter_coeff391_a(rf_filter_coeff391_a), 
    .rf_filter_coeff391_b(rf_filter_coeff391_b), 
    .rf_filter_coeff392_a(rf_filter_coeff392_a), 
    .rf_filter_coeff392_b(rf_filter_coeff392_b), 
    .rf_filter_coeff393_a(rf_filter_coeff393_a), 
    .rf_filter_coeff393_b(rf_filter_coeff393_b), 
    .rf_filter_coeff394_a(rf_filter_coeff394_a), 
    .rf_filter_coeff394_b(rf_filter_coeff394_b), 
    .rf_filter_coeff395_a(rf_filter_coeff395_a), 
    .rf_filter_coeff395_b(rf_filter_coeff395_b), 
    .rf_filter_coeff396_a(rf_filter_coeff396_a), 
    .rf_filter_coeff396_b(rf_filter_coeff396_b), 
    .rf_filter_coeff397_a(rf_filter_coeff397_a), 
    .rf_filter_coeff397_b(rf_filter_coeff397_b), 
    .rf_filter_coeff398_a(rf_filter_coeff398_a), 
    .rf_filter_coeff398_b(rf_filter_coeff398_b), 
    .rf_filter_coeff399_a(rf_filter_coeff399_a), 
    .rf_filter_coeff399_b(rf_filter_coeff399_b), 
    .rf_filter_coeff400_a(rf_filter_coeff400_a), 
    .rf_filter_coeff400_b(rf_filter_coeff400_b), 
    .rf_filter_coeff401_a(rf_filter_coeff401_a), 
    .rf_filter_coeff401_b(rf_filter_coeff401_b), 
    .rf_filter_coeff402_a(rf_filter_coeff402_a), 
    .rf_filter_coeff402_b(rf_filter_coeff402_b), 
    .rf_filter_coeff403_a(rf_filter_coeff403_a), 
    .rf_filter_coeff403_b(rf_filter_coeff403_b), 
    .rf_filter_coeff404_a(rf_filter_coeff404_a), 
    .rf_filter_coeff404_b(rf_filter_coeff404_b), 
    .rf_filter_coeff405_a(rf_filter_coeff405_a), 
    .rf_filter_coeff405_b(rf_filter_coeff405_b), 
    .rf_filter_coeff406_a(rf_filter_coeff406_a), 
    .rf_filter_coeff406_b(rf_filter_coeff406_b), 
    .rf_filter_coeff407_a(rf_filter_coeff407_a), 
    .rf_filter_coeff407_b(rf_filter_coeff407_b), 
    .rf_filter_coeff408_a(rf_filter_coeff408_a), 
    .rf_filter_coeff408_b(rf_filter_coeff408_b), 
    .rf_filter_coeff409_a(rf_filter_coeff409_a), 
    .rf_filter_coeff409_b(rf_filter_coeff409_b), 
    .rf_filter_coeff410_a(rf_filter_coeff410_a), 
    .rf_filter_coeff410_b(rf_filter_coeff410_b), 
    .rf_filter_coeff411_a(rf_filter_coeff411_a), 
    .rf_filter_coeff411_b(rf_filter_coeff411_b), 
    .rf_filter_coeff412_a(rf_filter_coeff412_a), 
    .rf_filter_coeff412_b(rf_filter_coeff412_b), 
    .rf_filter_coeff413_a(rf_filter_coeff413_a), 
    .rf_filter_coeff413_b(rf_filter_coeff413_b), 
    .rf_filter_coeff414_a(rf_filter_coeff414_a), 
    .rf_filter_coeff414_b(rf_filter_coeff414_b), 
    .rf_filter_coeff415_a(rf_filter_coeff415_a), 
    .rf_filter_coeff415_b(rf_filter_coeff415_b), 
    .rf_filter_coeff416_a(rf_filter_coeff416_a), 
    .rf_filter_coeff416_b(rf_filter_coeff416_b), 
    .rf_filter_coeff417_a(rf_filter_coeff417_a), 
    .rf_filter_coeff417_b(rf_filter_coeff417_b), 
    .rf_filter_coeff418_a(rf_filter_coeff418_a), 
    .rf_filter_coeff418_b(rf_filter_coeff418_b), 
    .rf_filter_coeff419_a(rf_filter_coeff419_a), 
    .rf_filter_coeff419_b(rf_filter_coeff419_b), 
    .rf_filter_coeff420_a(rf_filter_coeff420_a), 
    .rf_filter_coeff420_b(rf_filter_coeff420_b), 
    .rf_filter_coeff421_a(rf_filter_coeff421_a), 
    .rf_filter_coeff421_b(rf_filter_coeff421_b), 
    .rf_filter_coeff422_a(rf_filter_coeff422_a), 
    .rf_filter_coeff422_b(rf_filter_coeff422_b), 
    .rf_filter_coeff423_a(rf_filter_coeff423_a), 
    .rf_filter_coeff423_b(rf_filter_coeff423_b), 
    .rf_filter_coeff424_a(rf_filter_coeff424_a), 
    .rf_filter_coeff424_b(rf_filter_coeff424_b), 
    .rf_filter_coeff425_a(rf_filter_coeff425_a), 
    .rf_filter_coeff425_b(rf_filter_coeff425_b), 
    .rf_filter_coeff426_a(rf_filter_coeff426_a), 
    .rf_filter_coeff426_b(rf_filter_coeff426_b), 
    .rf_filter_coeff427_a(rf_filter_coeff427_a), 
    .rf_filter_coeff427_b(rf_filter_coeff427_b), 
    .rf_filter_coeff428_a(rf_filter_coeff428_a), 
    .rf_filter_coeff428_b(rf_filter_coeff428_b), 
    .rf_filter_coeff429_a(rf_filter_coeff429_a), 
    .rf_filter_coeff429_b(rf_filter_coeff429_b), 
    .rf_filter_coeff430_a(rf_filter_coeff430_a), 
    .rf_filter_coeff430_b(rf_filter_coeff430_b), 
    .rf_filter_coeff431_a(rf_filter_coeff431_a), 
    .rf_filter_coeff431_b(rf_filter_coeff431_b), 
    .rf_filter_coeff432_a(rf_filter_coeff432_a), 
    .rf_filter_coeff432_b(rf_filter_coeff432_b), 
    .rf_filter_coeff433_a(rf_filter_coeff433_a), 
    .rf_filter_coeff433_b(rf_filter_coeff433_b), 
    .rf_filter_coeff434_a(rf_filter_coeff434_a), 
    .rf_filter_coeff434_b(rf_filter_coeff434_b), 
    .rf_filter_coeff435_a(rf_filter_coeff435_a), 
    .rf_filter_coeff435_b(rf_filter_coeff435_b), 
    .rf_filter_coeff436_a(rf_filter_coeff436_a), 
    .rf_filter_coeff436_b(rf_filter_coeff436_b), 
    .rf_filter_coeff437_a(rf_filter_coeff437_a), 
    .rf_filter_coeff437_b(rf_filter_coeff437_b), 
    .rf_filter_coeff438_a(rf_filter_coeff438_a), 
    .rf_filter_coeff438_b(rf_filter_coeff438_b), 
    .rf_filter_coeff439_a(rf_filter_coeff439_a), 
    .rf_filter_coeff439_b(rf_filter_coeff439_b), 
    .rf_filter_coeff440_a(rf_filter_coeff440_a), 
    .rf_filter_coeff440_b(rf_filter_coeff440_b), 
    .rf_filter_coeff441_a(rf_filter_coeff441_a), 
    .rf_filter_coeff441_b(rf_filter_coeff441_b), 
    .rf_filter_coeff442_a(rf_filter_coeff442_a), 
    .rf_filter_coeff442_b(rf_filter_coeff442_b), 
    .rf_filter_coeff443_a(rf_filter_coeff443_a), 
    .rf_filter_coeff443_b(rf_filter_coeff443_b), 
    .rf_filter_coeff444_a(rf_filter_coeff444_a), 
    .rf_filter_coeff444_b(rf_filter_coeff444_b), 
    .rf_filter_coeff445_a(rf_filter_coeff445_a), 
    .rf_filter_coeff445_b(rf_filter_coeff445_b), 
    .rf_filter_coeff446_a(rf_filter_coeff446_a), 
    .rf_filter_coeff446_b(rf_filter_coeff446_b), 
    .rf_filter_coeff447_a(rf_filter_coeff447_a), 
    .rf_filter_coeff447_b(rf_filter_coeff447_b), 
    .rf_filter_coeff448_a(rf_filter_coeff448_a), 
    .rf_filter_coeff448_b(rf_filter_coeff448_b), 
    .rf_filter_coeff449_a(rf_filter_coeff449_a), 
    .rf_filter_coeff449_b(rf_filter_coeff449_b), 
    .rf_filter_coeff450_a(rf_filter_coeff450_a), 
    .rf_filter_coeff450_b(rf_filter_coeff450_b), 
    .rf_filter_coeff451_a(rf_filter_coeff451_a), 
    .rf_filter_coeff451_b(rf_filter_coeff451_b), 
    .rf_filter_coeff452_a(rf_filter_coeff452_a), 
    .rf_filter_coeff452_b(rf_filter_coeff452_b), 
    .rf_filter_coeff453_a(rf_filter_coeff453_a), 
    .rf_filter_coeff453_b(rf_filter_coeff453_b), 
    .rf_filter_coeff454_a(rf_filter_coeff454_a), 
    .rf_filter_coeff454_b(rf_filter_coeff454_b), 
    .rf_filter_coeff455_a(rf_filter_coeff455_a), 
    .rf_filter_coeff455_b(rf_filter_coeff455_b), 
    .rf_filter_coeff456_a(rf_filter_coeff456_a), 
    .rf_filter_coeff456_b(rf_filter_coeff456_b), 
    .rf_filter_coeff457_a(rf_filter_coeff457_a), 
    .rf_filter_coeff457_b(rf_filter_coeff457_b), 
    .rf_filter_coeff458_a(rf_filter_coeff458_a), 
    .rf_filter_coeff458_b(rf_filter_coeff458_b), 
    .rf_filter_coeff459_a(rf_filter_coeff459_a), 
    .rf_filter_coeff459_b(rf_filter_coeff459_b), 
    .rf_filter_coeff460_a(rf_filter_coeff460_a), 
    .rf_filter_coeff460_b(rf_filter_coeff460_b), 
    .rf_filter_coeff461_a(rf_filter_coeff461_a), 
    .rf_filter_coeff461_b(rf_filter_coeff461_b), 
    .rf_filter_coeff462_a(rf_filter_coeff462_a), 
    .rf_filter_coeff462_b(rf_filter_coeff462_b), 
    .rf_filter_coeff463_a(rf_filter_coeff463_a), 
    .rf_filter_coeff463_b(rf_filter_coeff463_b), 
    .rf_filter_coeff464_a(rf_filter_coeff464_a), 
    .rf_filter_coeff464_b(rf_filter_coeff464_b), 
    .rf_filter_coeff465_a(rf_filter_coeff465_a), 
    .rf_filter_coeff465_b(rf_filter_coeff465_b), 
    .rf_filter_coeff466_a(rf_filter_coeff466_a), 
    .rf_filter_coeff466_b(rf_filter_coeff466_b), 
    .rf_filter_coeff467_a(rf_filter_coeff467_a), 
    .rf_filter_coeff467_b(rf_filter_coeff467_b), 
    .rf_filter_coeff468_a(rf_filter_coeff468_a), 
    .rf_filter_coeff468_b(rf_filter_coeff468_b), 
    .rf_filter_coeff469_a(rf_filter_coeff469_a), 
    .rf_filter_coeff469_b(rf_filter_coeff469_b), 
    .rf_filter_coeff470_a(rf_filter_coeff470_a), 
    .rf_filter_coeff470_b(rf_filter_coeff470_b), 
    .rf_filter_coeff471_a(rf_filter_coeff471_a), 
    .rf_filter_coeff471_b(rf_filter_coeff471_b), 
    .rf_filter_coeff472_a(rf_filter_coeff472_a), 
    .rf_filter_coeff472_b(rf_filter_coeff472_b), 
    .rf_filter_coeff473_a(rf_filter_coeff473_a), 
    .rf_filter_coeff473_b(rf_filter_coeff473_b), 
    .rf_filter_coeff474_a(rf_filter_coeff474_a), 
    .rf_filter_coeff474_b(rf_filter_coeff474_b), 
    .rf_filter_coeff475_a(rf_filter_coeff475_a), 
    .rf_filter_coeff475_b(rf_filter_coeff475_b), 
    .rf_filter_coeff476_a(rf_filter_coeff476_a), 
    .rf_filter_coeff476_b(rf_filter_coeff476_b), 
    .rf_filter_coeff477_a(rf_filter_coeff477_a), 
    .rf_filter_coeff477_b(rf_filter_coeff477_b), 
    .rf_filter_coeff478_a(rf_filter_coeff478_a), 
    .rf_filter_coeff478_b(rf_filter_coeff478_b), 
    .rf_filter_coeff479_a(rf_filter_coeff479_a), 
    .rf_filter_coeff479_b(rf_filter_coeff479_b), 
    .rf_filter_coeff480_a(rf_filter_coeff480_a), 
    .rf_filter_coeff480_b(rf_filter_coeff480_b), 
    .rf_filter_coeff481_a(rf_filter_coeff481_a), 
    .rf_filter_coeff481_b(rf_filter_coeff481_b), 
    .rf_filter_coeff482_a(rf_filter_coeff482_a), 
    .rf_filter_coeff482_b(rf_filter_coeff482_b), 
    .rf_filter_coeff483_a(rf_filter_coeff483_a), 
    .rf_filter_coeff483_b(rf_filter_coeff483_b), 
    .rf_filter_coeff484_a(rf_filter_coeff484_a), 
    .rf_filter_coeff484_b(rf_filter_coeff484_b), 
    .rf_filter_coeff485_a(rf_filter_coeff485_a), 
    .rf_filter_coeff485_b(rf_filter_coeff485_b), 
    .rf_filter_coeff486_a(rf_filter_coeff486_a), 
    .rf_filter_coeff486_b(rf_filter_coeff486_b), 
    .rf_filter_coeff487_a(rf_filter_coeff487_a), 
    .rf_filter_coeff487_b(rf_filter_coeff487_b), 
    .rf_filter_coeff488_a(rf_filter_coeff488_a), 
    .rf_filter_coeff488_b(rf_filter_coeff488_b), 
    .rf_filter_coeff489_a(rf_filter_coeff489_a), 
    .rf_filter_coeff489_b(rf_filter_coeff489_b), 
    .rf_filter_coeff490_a(rf_filter_coeff490_a), 
    .rf_filter_coeff490_b(rf_filter_coeff490_b), 
    .rf_filter_coeff491_a(rf_filter_coeff491_a), 
    .rf_filter_coeff491_b(rf_filter_coeff491_b), 
    .rf_filter_coeff492_a(rf_filter_coeff492_a), 
    .rf_filter_coeff492_b(rf_filter_coeff492_b), 
    .rf_filter_coeff493_a(rf_filter_coeff493_a), 
    .rf_filter_coeff493_b(rf_filter_coeff493_b), 
    .rf_filter_coeff494_a(rf_filter_coeff494_a), 
    .rf_filter_coeff494_b(rf_filter_coeff494_b), 
    .rf_filter_coeff495_a(rf_filter_coeff495_a), 
    .rf_filter_coeff495_b(rf_filter_coeff495_b), 
    .rf_filter_coeff496_a(rf_filter_coeff496_a), 
    .rf_filter_coeff496_b(rf_filter_coeff496_b), 
    .rf_filter_coeff497_a(rf_filter_coeff497_a), 
    .rf_filter_coeff497_b(rf_filter_coeff497_b), 
    .rf_filter_coeff498_a(rf_filter_coeff498_a), 
    .rf_filter_coeff498_b(rf_filter_coeff498_b), 
    .rf_filter_coeff499_a(rf_filter_coeff499_a), 
    .rf_filter_coeff499_b(rf_filter_coeff499_b), 
    .rf_filter_coeff500_a(rf_filter_coeff500_a), 
    .rf_filter_coeff500_b(rf_filter_coeff500_b), 
    .rf_filter_coeff501_a(rf_filter_coeff501_a), 
    .rf_filter_coeff501_b(rf_filter_coeff501_b), 
    .rf_filter_coeff502_a(rf_filter_coeff502_a), 
    .rf_filter_coeff502_b(rf_filter_coeff502_b), 
    .rf_filter_coeff503_a(rf_filter_coeff503_a), 
    .rf_filter_coeff503_b(rf_filter_coeff503_b), 
    .rf_filter_coeff504_a(rf_filter_coeff504_a), 
    .rf_filter_coeff504_b(rf_filter_coeff504_b), 
    .rf_filter_coeff505_a(rf_filter_coeff505_a), 
    .rf_filter_coeff505_b(rf_filter_coeff505_b), 
    .rf_filter_coeff506_a(rf_filter_coeff506_a), 
    .rf_filter_coeff506_b(rf_filter_coeff506_b), 
    .rf_filter_coeff507_a(rf_filter_coeff507_a), 
    .rf_filter_coeff507_b(rf_filter_coeff507_b), 
    .rf_filter_coeff508_a(rf_filter_coeff508_a), 
    .rf_filter_coeff508_b(rf_filter_coeff508_b), 
    .rf_filter_coeff509_a(rf_filter_coeff509_a), 
    .rf_filter_coeff509_b(rf_filter_coeff509_b), 
    .rf_filter_coeff510_a(rf_filter_coeff510_a), 
    .rf_filter_coeff510_b(rf_filter_coeff510_b), 
    .rf_filter_coeff511_a(rf_filter_coeff511_a), 
    .rf_filter_coeff511_b(rf_filter_coeff511_b)
    );
//***********************************************************************************


endmodule
