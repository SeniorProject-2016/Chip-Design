`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    12:59:12 06/06/2015 
// Design Name: 
// Module Name:    register 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module register(
    input clk,
    input rst,
    input op,
    input [9:0] addr,
    input [31:0] wdata,
    input rts,
    output rtr,
    output [31:0] rdata,
    output xfc,
    input i2s_overrun
    );


endmodule
