//////////////////////////////////////////////////////////////////////////////////
// Module Name:             filter_storage.v
// Create Date:             ??? 
// Last Modification:       3/25/2016
// Author:                  Dhruvit Naik
// Description:             ????
//////////////////////////////////////////////////////////////////////////////////

`timescale 1ns / 1ps

module filter_storage( clk, rst_n, wren, wrptr, wrdata, rden, rdptr, rddata
    );

    input								    clk;
    input								    rst_n;
    input								    wren;
    input		    [8:0]					wrptr;
    input		    [31:0]				    wrdata;
    input								    rden;
    input		    [8:0]					rdptr;
    output	        [31:0]				    rddata;

    localparam	                            DEPTH = 511; //2^9 <= 16'b0; 512
    localparam	                            WIDTH = 31; 

    reg	            [WIDTH:0]               ram [DEPTH:0];
    reg	            [WIDTH:0]               rddata;	


    always @(posedge clk or negedge rst_n)
    begin
        if (!rst_n)
        begin
             ram[0] <= 16'b0;
             ram[1] <= 16'b0; 
             ram[2] <= 16'b0; 
             ram[3] <= 16'b0;  
             ram[4] <= 16'b0; 
             ram[5] <= 16'b0; 
             ram[6] <= 16'b0; 
             ram[7] <= 16'b0; 
             ram[8] <= 16'b0;  
             ram[9] <= 16'b0;
             ram[10] <= 16'b0; 
             ram[11] <= 16'b0; 
             ram[12] <= 16'b0;  
             ram[13] <= 16'b0;  
             ram[14] <= 16'b0; 
             ram[15] <= 16'b0; 
             ram[16] <= 16'b0; 
             ram[17] <= 16'b0;  
             ram[18] <= 16'b0; 
             ram[19] <= 16'b0;
             ram[20] <= 16'b0; 
             ram[21] <= 16'b0; 
             ram[22] <= 16'b0; 
             ram[23] <= 16'b0; 
             ram[24] <= 16'b0; 
             ram[25] <= 16'b0; 
             ram[26] <= 16'b0; 
             ram[27] <= 16'b0; 
             ram[28] <= 16'b0; 
             ram[29] <= 16'b0; 
             ram[30] <= 16'b0; 
             ram[31] <= 16'b0; 
             ram[32] <= 16'b0; 
             ram[33] <= 16'b0; 
             ram[34] <= 16'b0; 
             ram[35] <= 16'b0; 
             ram[36] <= 16'b0; 
             ram[37] <= 16'b0; 
             ram[38] <= 16'b0; 
             ram[39] <= 16'b0; 
             ram[40] <= 16'b0; 
             ram[41] <= 16'b0; 
             ram[42] <= 16'b0; 
             ram[43] <= 16'b0; 
             ram[44] <= 16'b0; 
             ram[45] <= 16'b0; 
             ram[46] <= 16'b0; 
             ram[47] <= 16'b0; 
             ram[48] <= 16'b0; 
             ram[49] <= 16'b0; 
             ram[50] <= 16'b0; 
             ram[51] <= 16'b0; 
             ram[52] <= 16'b0; 
             ram[53] <= 16'b0; 
             ram[54] <= 16'b0; 
             ram[55] <= 16'b0; 
             ram[56] <= 16'b0; 
             ram[57] <= 16'b0; 
             ram[58] <= 16'b0; 
             ram[59] <= 16'b0; 
             ram[60] <= 16'b0; 
             ram[61] <= 16'b0; 
             ram[62] <= 16'b0; 
             ram[63] <= 16'b0; 
             ram[64] <= 16'b0; 
             ram[65] <= 16'b0; 
             ram[66] <= 16'b0; 
             ram[67] <= 16'b0; 
             ram[68] <= 16'b0; 
             ram[69] <= 16'b0; 
             ram[70] <= 16'b0; 
             ram[71] <= 16'b0; 
             ram[72] <= 16'b0; 
             ram[73] <= 16'b0; 
             ram[74] <= 16'b0; 
             ram[75] <= 16'b0; 
             ram[76] <= 16'b0; 
             ram[77] <= 16'b0; 
             ram[78] <= 16'b0; 
             ram[79] <= 16'b0; 
             ram[80] <= 16'b0; 
             ram[81] <= 16'b0; 
             ram[82] <= 16'b0; 
             ram[83] <= 16'b0; 
             ram[84] <= 16'b0; 
             ram[85] <= 16'b0; 
             ram[86] <= 16'b0; 
             ram[87] <= 16'b0; 
             ram[88] <= 16'b0; 
             ram[89] <= 16'b0; 
             ram[90] <= 16'b0; 
             ram[91] <= 16'b0; 
             ram[92] <= 16'b0; 
             ram[93] <= 16'b0; 
             ram[94] <= 16'b0; 
             ram[95] <= 16'b0; 
             ram[96] <= 16'b0; 
             ram[97] <= 16'b0; 
             ram[98] <= 16'b0; 
             ram[99] <= 16'b0; 
             ram[100] <= 16'b0;
             ram[101] <= 16'b0; 
             ram[102] <= 16'b0; 
             ram[103] <= 16'b0; 
             ram[104] <= 16'b0; 
             ram[105] <= 16'b0; 
             ram[106] <= 16'b0; 
             ram[107] <= 16'b0; 
             ram[108] <= 16'b0; 
             ram[109] <= 16'b0; 
             ram[110] <= 16'b0; 
             ram[111] <= 16'b0; 
             ram[112] <= 16'b0; 
             ram[113] <= 16'b0; 
             ram[114] <= 16'b0; 
             ram[115] <= 16'b0; 
             ram[116] <= 16'b0; 
             ram[117] <= 16'b0; 
             ram[118] <= 16'b0; 
             ram[119] <= 16'b0; 
             ram[120] <= 16'b0; 
             ram[121] <= 16'b0; 
             ram[122] <= 16'b0; 
             ram[123] <= 16'b0; 
             ram[124] <= 16'b0; 
             ram[125] <= 16'b0; 
             ram[126] <= 16'b0; 
             ram[127] <= 16'b0; 
             ram[128] <= 16'b0; 
             ram[129] <= 16'b0; 
             ram[130] <= 16'b0; 
             ram[131] <= 16'b0; 
             ram[132] <= 16'b0; 
             ram[133] <= 16'b0; 
             ram[134] <= 16'b0; 
             ram[135] <= 16'b0; 
             ram[136] <= 16'b0; 
             ram[137] <= 16'b0; 
             ram[138] <= 16'b0; 
             ram[139] <= 16'b0; 
             ram[140] <= 16'b0; 
             ram[141] <= 16'b0; 
             ram[142] <= 16'b0; 
             ram[143] <= 16'b0; 
             ram[144] <= 16'b0; 
             ram[145] <= 16'b0; 
             ram[146] <= 16'b0; 
             ram[147] <= 16'b0; 
             ram[148] <= 16'b0; 
             ram[149] <= 16'b0; 
             ram[150] <= 16'b0; 
             ram[151] <= 16'b0; 
             ram[152] <= 16'b0; 
             ram[153] <= 16'b0; 
             ram[154] <= 16'b0; 
             ram[155] <= 16'b0; 
             ram[156] <= 16'b0; 
             ram[157] <= 16'b0; 
             ram[158] <= 16'b0; 
             ram[159] <= 16'b0; 
             ram[160] <= 16'b0; 
             ram[161] <= 16'b0; 
             ram[162] <= 16'b0; 
             ram[163] <= 16'b0; 
             ram[164] <= 16'b0; 
             ram[165] <= 16'b0; 
             ram[166] <= 16'b0; 
             ram[167] <= 16'b0; 
             ram[168] <= 16'b0; 
             ram[169] <= 16'b0; 
             ram[170] <= 16'b0; 
             ram[171] <= 16'b0; 
             ram[172] <= 16'b0; 
             ram[173] <= 16'b0; 
             ram[174] <= 16'b0; 
             ram[175] <= 16'b0; 
             ram[176] <= 16'b0; 
             ram[177] <= 16'b0; 
             ram[178] <= 16'b0; 
             ram[179] <= 16'b0; 
             ram[180] <= 16'b0; 
             ram[181] <= 16'b0; 
             ram[182] <= 16'b0; 
             ram[183] <= 16'b0; 
             ram[184] <= 16'b0; 
             ram[185] <= 16'b0; 
             ram[186] <= 16'b0; 
             ram[187] <= 16'b0; 
             ram[188] <= 16'b0; 
             ram[189] <= 16'b0; 
             ram[190] <= 16'b0; 
             ram[191] <= 16'b0; 
             ram[192] <= 16'b0; 
             ram[193] <= 16'b0; 
             ram[194] <= 16'b0; 
             ram[195] <= 16'b0; 
             ram[196] <= 16'b0; 
             ram[197] <= 16'b0; 
             ram[198] <= 16'b0; 
             ram[199] <= 16'b0; 
             ram[200] <= 16'b0; 
             ram[201] <= 16'b0; 
             ram[202] <= 16'b0; 
             ram[203] <= 16'b0; 
             ram[204] <= 16'b0; 
             ram[205] <= 16'b0; 
             ram[206] <= 16'b0; 
             ram[207] <= 16'b0; 
             ram[208] <= 16'b0; 
             ram[209] <= 16'b0; 
             ram[210] <= 16'b0; 
             ram[211] <= 16'b0; 
             ram[212] <= 16'b0; 
             ram[213] <= 16'b0; 
             ram[214] <= 16'b0; 
             ram[215] <= 16'b0; 
             ram[216] <= 16'b0; 
             ram[217] <= 16'b0; 
             ram[218] <= 16'b0; 
             ram[219] <= 16'b0; 
             ram[220] <= 16'b0; 
             ram[221] <= 16'b0; 
             ram[222] <= 16'b0; 
             ram[223] <= 16'b0; 
             ram[224] <= 16'b0; 
             ram[225] <= 16'b0; 
             ram[226] <= 16'b0; 
             ram[227] <= 16'b0; 
             ram[228] <= 16'b0; 
             ram[229] <= 16'b0; 
             ram[230] <= 16'b0; 
             ram[231] <= 16'b0; 
             ram[232] <= 16'b0; 
             ram[233] <= 16'b0; 
             ram[234] <= 16'b0; 
             ram[235] <= 16'b0; 
             ram[236] <= 16'b0; 
             ram[237] <= 16'b0; 
             ram[238] <= 16'b0; 
             ram[239] <= 16'b0; 
             ram[240] <= 16'b0; 
             ram[241] <= 16'b0; 
             ram[242] <= 16'b0; 
             ram[243] <= 16'b0; 
             ram[244] <= 16'b0; 
             ram[245] <= 16'b0; 
             ram[246] <= 16'b0; 
             ram[247] <= 16'b0; 
             ram[248] <= 16'b0; 
             ram[249] <= 16'b0; 
             ram[250] <= 16'b0; 
             ram[251] <= 16'b0; 
             ram[252] <= 16'b0; 
             ram[253] <= 16'b0; 
             ram[254] <= 16'b0; 
             ram[255] <= 16'b0; 
             ram[256] <= 16'b0; 
             ram[257] <= 16'b0; 
             ram[258] <= 16'b0; 
             ram[259] <= 16'b0; 
             ram[260] <= 16'b0; 
             ram[261] <= 16'b0; 
             ram[262] <= 16'b0; 
             ram[263] <= 16'b0; 
             ram[264] <= 16'b0; 
             ram[265] <= 16'b0; 
             ram[266] <= 16'b0; 
             ram[267] <= 16'b0; 
             ram[268] <= 16'b0; 
             ram[269] <= 16'b0; 
             ram[270] <= 16'b0; 
             ram[271] <= 16'b0; 
             ram[272] <= 16'b0; 
             ram[273] <= 16'b0; 
             ram[274] <= 16'b0; 
             ram[275] <= 16'b0; 
             ram[276] <= 16'b0; 
             ram[277] <= 16'b0; 
             ram[278] <= 16'b0; 
             ram[279] <= 16'b0; 
             ram[280] <= 16'b0; 
             ram[281] <= 16'b0; 
             ram[282] <= 16'b0; 
             ram[283] <= 16'b0; 
             ram[284] <= 16'b0; 
             ram[285] <= 16'b0; 
             ram[286] <= 16'b0; 
             ram[287] <= 16'b0; 
             ram[288] <= 16'b0; 
             ram[289] <= 16'b0; 
             ram[290] <= 16'b0; 
             ram[291] <= 16'b0; 
             ram[292] <= 16'b0; 
             ram[293] <= 16'b0; 
             ram[294] <= 16'b0; 
             ram[295] <= 16'b0; 
             ram[296] <= 16'b0; 
             ram[297] <= 16'b0; 
             ram[298] <= 16'b0; 
             ram[299] <= 16'b0; 
             ram[300] <= 16'b0; 
             ram[301] <= 16'b0; 
             ram[302] <= 16'b0; 
             ram[303] <= 16'b0; 
             ram[304] <= 16'b0; 
             ram[305] <= 16'b0; 
             ram[306] <= 16'b0; 
             ram[307] <= 16'b0; 
             ram[308] <= 16'b0; 
             ram[309] <= 16'b0; 
             ram[310] <= 16'b0; 
             ram[311] <= 16'b0; 
             ram[312] <= 16'b0; 
             ram[313] <= 16'b0; 
             ram[314] <= 16'b0; 
             ram[315] <= 16'b0; 
             ram[316] <= 16'b0; 
             ram[317] <= 16'b0; 
             ram[318] <= 16'b0; 
             ram[319] <= 16'b0; 
             ram[320] <= 16'b0; 
             ram[321] <= 16'b0; 
             ram[322] <= 16'b0; 
             ram[323] <= 16'b0; 
             ram[324] <= 16'b0; 
             ram[325] <= 16'b0; 
             ram[326] <= 16'b0; 
             ram[327] <= 16'b0; 
             ram[328] <= 16'b0; 
             ram[329] <= 16'b0; 
             ram[330] <= 16'b0; 
             ram[331] <= 16'b0; 
             ram[332] <= 16'b0; 
             ram[333] <= 16'b0; 
             ram[334] <= 16'b0; 
             ram[335] <= 16'b0; 
             ram[336] <= 16'b0; 
             ram[337] <= 16'b0; 
             ram[338] <= 16'b0; 
             ram[339] <= 16'b0; 
             ram[340] <= 16'b0; 
             ram[341] <= 16'b0; 
             ram[342] <= 16'b0; 
             ram[343] <= 16'b0; 
             ram[344] <= 16'b0; 
             ram[345] <= 16'b0; 
             ram[346] <= 16'b0; 
             ram[347] <= 16'b0; 
             ram[348] <= 16'b0; 
             ram[349] <= 16'b0; 
             ram[350] <= 16'b0; 
             ram[351] <= 16'b0; 
             ram[352] <= 16'b0; 
             ram[353] <= 16'b0; 
             ram[354] <= 16'b0; 
             ram[355] <= 16'b0; 
             ram[356] <= 16'b0; 
             ram[357] <= 16'b0; 
             ram[358] <= 16'b0; 
             ram[359] <= 16'b0; 
             ram[360] <= 16'b0; 
             ram[361] <= 16'b0; 
             ram[362] <= 16'b0; 
             ram[363] <= 16'b0; 
             ram[364] <= 16'b0; 
             ram[365] <= 16'b0; 
             ram[366] <= 16'b0; 
             ram[367] <= 16'b0; 
             ram[368] <= 16'b0; 
             ram[369] <= 16'b0; 
             ram[370] <= 16'b0; 
             ram[371] <= 16'b0; 
             ram[372] <= 16'b0; 
             ram[373] <= 16'b0; 
             ram[374] <= 16'b0; 
             ram[375] <= 16'b0; 
             ram[376] <= 16'b0; 
             ram[377] <= 16'b0; 
             ram[378] <= 16'b0; 
             ram[379] <= 16'b0; 
             ram[380] <= 16'b0; 
             ram[381] <= 16'b0; 
             ram[382] <= 16'b0; 
             ram[383] <= 16'b0; 
             ram[384] <= 16'b0; 
             ram[385] <= 16'b0; 
             ram[386] <= 16'b0; 
             ram[387] <= 16'b0; 
             ram[388] <= 16'b0; 
             ram[389] <= 16'b0; 
             ram[390] <= 16'b0; 
             ram[391] <= 16'b0; 
             ram[392] <= 16'b0; 
             ram[393] <= 16'b0; 
             ram[394] <= 16'b0; 
             ram[395] <= 16'b0; 
             ram[396] <= 16'b0; 
             ram[397] <= 16'b0; 
             ram[398] <= 16'b0; 
             ram[399] <= 16'b0; 
             ram[400] <= 16'b0; 
             ram[401] <= 16'b0; 
             ram[402] <= 16'b0; 
             ram[403] <= 16'b0; 
             ram[404] <= 16'b0; 
             ram[405] <= 16'b0; 
             ram[406] <= 16'b0; 
             ram[407] <= 16'b0; 
             ram[408] <= 16'b0; 
             ram[409] <= 16'b0; 
             ram[410] <= 16'b0; 
             ram[411] <= 16'b0; 
             ram[412] <= 16'b0; 
             ram[413] <= 16'b0; 
             ram[414] <= 16'b0; 
             ram[415] <= 16'b0; 
             ram[416] <= 16'b0; 
             ram[417] <= 16'b0; 
             ram[418] <= 16'b0; 
             ram[419] <= 16'b0; 
             ram[420] <= 16'b0; 
             ram[421] <= 16'b0; 
             ram[422] <= 16'b0; 
             ram[423] <= 16'b0; 
             ram[424] <= 16'b0; 
             ram[425] <= 16'b0; 
             ram[426] <= 16'b0; 
             ram[427] <= 16'b0; 
             ram[428] <= 16'b0; 
             ram[429] <= 16'b0; 
             ram[430] <= 16'b0; 
             ram[431] <= 16'b0; 
             ram[432] <= 16'b0; 
             ram[433] <= 16'b0; 
             ram[434] <= 16'b0; 
             ram[435] <= 16'b0; 
             ram[436] <= 16'b0; 
             ram[437] <= 16'b0; 
             ram[438] <= 16'b0; 
             ram[439] <= 16'b0; 
             ram[440] <= 16'b0; 
             ram[441] <= 16'b0; 
             ram[442] <= 16'b0; 
             ram[443] <= 16'b0; 
             ram[444] <= 16'b0; 
             ram[445] <= 16'b0; 
             ram[446] <= 16'b0; 
             ram[447] <= 16'b0; 
             ram[448] <= 16'b0; 
             ram[449] <= 16'b0; 
             ram[450] <= 16'b0; 
             ram[451] <= 16'b0; 
             ram[452] <= 16'b0; 
             ram[453] <= 16'b0; 
             ram[454] <= 16'b0; 
             ram[455] <= 16'b0; 
             ram[456] <= 16'b0; 
             ram[457] <= 16'b0; 
             ram[458] <= 16'b0; 
             ram[459] <= 16'b0; 
             ram[460] <= 16'b0; 
             ram[461] <= 16'b0; 
             ram[462] <= 16'b0; 
             ram[463] <= 16'b0; 
             ram[464] <= 16'b0; 
             ram[465] <= 16'b0; 
             ram[466] <= 16'b0; 
             ram[467] <= 16'b0; 
             ram[468] <= 16'b0; 
             ram[469] <= 16'b0; 
             ram[470] <= 16'b0; 
             ram[471] <= 16'b0; 
             ram[472] <= 16'b0; 
             ram[473] <= 16'b0; 
             ram[474] <= 16'b0; 
             ram[475] <= 16'b0; 
             ram[476] <= 16'b0; 
             ram[477] <= 16'b0; 
             ram[478] <= 16'b0; 
             ram[479] <= 16'b0; 
             ram[480] <= 16'b0; 
             ram[481] <= 16'b0; 
             ram[482] <= 16'b0; 
             ram[483] <= 16'b0; 
             ram[484] <= 16'b0; 
             ram[485] <= 16'b0; 
             ram[486] <= 16'b0; 
             ram[487] <= 16'b0; 
             ram[488] <= 16'b0; 
             ram[489] <= 16'b0; 
             ram[490] <= 16'b0; 
             ram[491] <= 16'b0; 
             ram[492] <= 16'b0; 
             ram[493] <= 16'b0; 
             ram[494] <= 16'b0; 
             ram[495] <= 16'b0; 
             ram[496] <= 16'b0; 
             ram[497] <= 16'b0; 
             ram[498] <= 16'b0; 
             ram[499] <= 16'b0; 
             ram[500] <= 16'b0; 
             ram[501] <= 16'b0; 
             ram[502] <= 16'b0; 
             ram[503] <= 16'b0; 
             ram[504] <= 16'b0; 
             ram[505] <= 16'b0; 
             ram[506] <= 16'b0; 
             ram[507] <= 16'b0; 
             ram[508] <= 16'b0; 
             ram[509] <= 16'b0; 
             ram[510] <= 16'b0; 
             ram[511] <= 16'b0; 	
        end
        
        else if(wren)
            ram[wrptr] <= wrdata;

    end
        
    always @(posedge clk)
    begin
        if(rden)
            rddata <= ram[rdptr];
    end
        
endmodule
